��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�[� ��P4Xi�%�T��x�Y�c���ۣŤ�LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނf�Ey��ܷ��c�:o^L����@qґ��Jӣ.�
tٻС���7e�4{ȅ���8��R�FK�WQ_�i!�����o7�wby��<EK�)��S��{�Z-� q��6g"I��U=�p;��W�\H��P�S%�� ��YD- 8�bl�둄�=�1�E�b�B	�hWn���)Z�߄� ?�˺�>��p00꠷�����wŸE�x�E����*�<5���N5�P������=:�V�&z���ko։̿�#t΄�iЀkŶ�h�!!�h}�����S�@��q*��}m��1Cܖ����fT+(�x���>g�� 6�+��F�YS̢�~Dܞ}L[bu�a�P\�;�E^��33++�5�s�]y��M�_���8�:S�TQ09������:U���ꃅ�Y���
���S�-!`9���.z�������`�uŨUC�$]/W��ͮ��4|��/
��⭓r�X�������3_ͩ��}Ckll9Y�HMc?�?c��;�aJJ�"B��1L���8L�c���G��Q�FE��G��%2�l��`q�e�hʫ�-�O)�1�5"Hj���.4݂�����vlX����Hh@�zo��COz�ǚ���n�p�*Y dL�u�ϙ8@`���;�56n�ĥ]����C��t�n�-�����T-c^};Ycx1��ܳ�6���nŭ��ǋ�t9�h���>3b����uuO��k���"LP���;�ێ�H@ �}�����#�Tƽ̅��A����ܭu<��%ӵ�ci��^@̃Յ���N�cMW@��Pa��� W H-a~�i�Z�]KΎt<iOנ&�x�
_�F69��KF����L�75.�]�H��^�a�\nu���A�]";���Ϫ���A�"�Ep��} [���P�@���f�u�i�eD��7��²;T�K~����n�|�Į1&H���ލ�Td?��Iբo����y��w�k8@��*Nʵ�N���e'ҫ)C�5��b?���Gbd���m����?֫6[���a�G�NU�s�aK�zY+3ld&��$��^s*2�����<�TJ��H��]�G�]ӊ�%��6�N�B �'/`����2�����8�hI�(�@��͡�5���UfI!��є���ߔYݕub����g��E_�7��%tz���w��hl�qi��H�������5�im�w �j�-<"k�@�����D�%ǵt��������ʫ|Xy
�C@zu�2�o��\h�0p�^����IA�t7v,/h�h����&�� q(�7H\�VH<l��=��De6�P"��Q{�w�)� ��&���z�҆�ÑR��l �[�U�u,�OCx��铤���*�MCLa�ۭ��.����Xz���ߋCC%�}q/�q��0�B�^x��GW�3{��c*���_�Z���SBґ�؅J�@�C�O"�Q���Խ���%�۫���`�凣��k�X��iC������O~� R���l��V]S_�~��r@WR��9�S]����#�rpm5�J3�X�Q�G4������"���l}��3&JKlE#E�F$Y ����V
�V�p�6��K��n�#�a���М_
�B)W�fP;h�2s��\�[�Gq�呴�^�n�]�P��Hj��Z�}Q{[k�O�AΝOfr�mG!�ą,��A�v�FO�(�#�s�N��,?�IkA>��S�#�������q�-Szp� 	Mrg����q�[�1Q}�,R�Ѱ91�xb��.�=n7SQ8Qb��[��#���ZS��o�Q`��ף8�ʨ.�"�MFR�0��/���J�;�*�c'�2��aw5���@{;ۃ��Pzv�M�����#3(��u���Y�K�&�Gk�����-���MXUI��!�E������[ni����݉u��4��� 0X�8�Wob4�/�%��7?�_�h�~�y>��������D���oHn������Â��|-����)�E��[���{���`oGU�P��~�i�x���<�V)`�Һ���2��6��ւ�}б���o��ư��� ��2+mV�����^?�S��y�:(�СN|i��Q?��	w�~W���sI$R��?i�8�d��>,�	�~HŻI|���9�}Kԛ��@Pʅ"�}_*Zt���������'��Am�)��ЧKa$���e�#�a=[�ƺk#���L}m�*Afs�N���1��X��[���iyo�`U�ҕ�m��]��^`�z�g����5���i8"�8pSJ!�V��&�)�X��L*�u	ĵ���-�n=>�:�&��Sm�Jki>[;/�ʦ���/A���,`��- ]$�8f�>��TR��b�6��aҲ�6VȃJ������w.��
h�dSO\�Eƴ�Ƙ�w�P����� (0S��#EW�;���|}��¾r~7��ZQ�ݏ�l�'m��5�Wջ��큽�*l�x��k���j��V�\��3��إ��,{�2nA��\��,^�)q�5�+��j$|�I�F�D��ה��qdIy���
,4n�����6�펯 ������7o��Y���'<�|*�=M��:DJ{<b�x�k�8*���#ǌ����-A�e��{��Ԥ]/u��Z	8T�P�<��t}��������1x���>y��Z��J��-�J�l��R�\7���YS�+,�M�0�R>�ה�\�ms{��_�"�֥�	�L��k��D�;�G�mSL��[���^?�oβ,˜zr�B�tq�:&�l���N�/S[��2y/�����Ѹ�#�p<���D�dV@�̭ &}�GC��T�=1����>� {�����%�X#p����iU*�e��cE���'Y�NSc��0����$��E��*H��8���7=��&�G�G.�/����Զc�g#�k��?f�>yt7X�7�4�{��7�0�D^��E�T�V}��0��6�\����� ײ�ë��|��#��>�n�qn��??U�kD9Վq�I2 �9Ǉ���d�ߣ��YX1eLmm.��ح=·�P`����xY�+@��[���c��b�L	�9D�ȳ�s
o>�֯ܿ
º}/s<�G��� ��À���h~�s����'�t4Q���J��I�G��)��!5JÃ��I�u�M��[�o�/�.7�"�+`��ϔ�c�����������$��4�ZY��Z���Ph
��OԻ[kF�H~.��X�L�3��V�'t]M�0���8.��]?��

|���Ŷ����Qbw��x�dBQ��/e@M��O}B�/��*�ar!a��?�JMq?�*2���w��@2S�wq�f,N�0Z2�mZ��Zf��ʏ��	�6��'�L��eҳ��#���s��,ѸQ�����Lu�}!�~��Ȧ���+s�8��޼
�w�-���N���'_D#��h[�GD��m���h�Ĺ��-�Q��M�Ȑ�.fOfx�^�+�jw(2*�9�T膠���1>EFC���\,�� p)�����]�[�Z����G����i��DW�?��7)��i��p����0�Fd�GM��e���̳���#�O�R����Ūg��g�ƭ��@Æ���44���nTf���aw �+"���|l��$C����|+���.�-|ӹz�b.���_fY�jnU�iU�W�;rW�f��y��_�:�V�Qٯ�.0������[��<��X�a������!����דսw,�_�
�@�U��� �R�b嘩T� ���Gz�nx�K�P��wi�D����X��♭?Y����jʤ��gxEC\���/����P2�
^�&�����MU�A&/����Vpm����΀��_\$�����6H]՘1��
/����Q��L�B����Fu��1��[�01W�<�VW|!h�5��"���/ #_����e2�������8N�"^��@5lHN��yA��F�0Wv��� ��H�4�6kN*B/9���kJ(Y�8-��B�5�����2 �O$���I�W�}Q�Cq�|��q�t��v*Ț���Ԥ�M�Ɵ��SCs�ҙDY��?|"V��}��Y�BH�t��\���	i�A�q�厺d-� �v��P&+H>�N:����0��~�7�z��G� �.#��h��7���������]c�gR���E%����R�I,�>��!���Q��l��k�$�@�X@O&,��~]0��Ll;w+Ѻxп��F�>̄���}�+i��(�����;��zt��&��1�D����k�j̩W��	��TQU���!�T�)�Z�N�`4Y�9]�7J3�Eӟ�?�6NN�G��O���x��?�������p����d~5ca�¸��֪ȃ�FЄW˾������&U�a� r��J�}�,���
$0?����.��}4w2��#03�9o4���6�L6���$s�`�|���Z�8Â�����տmv�	<�M��A���Y�)b���e�5���?��l����8���w�sp��0Y�dP�ܔ�m�lƇ��.e�N����Z��B�3L�&˟�3΀A:A��m\P�
BL�"�@�J��E��C� ;U��ZI��)�zO��9�J�;�H͐8&&�z������J�N� )�B��?�%�k��k�WXc��C��!|Mlٌ�e�=W,����)j�.s؊�\04�q��e����c�a5;l8_`�  E4P��|jȲ���+���$j_�8�{~"�.!�����_��!��wκ�DcdI��f�f���"{�=���c(��C�� �d%}5�A�k
���D���͇�N.�!�g�;��<�}�$��a��HIH2��0țU��띌�J�,��:�:�"��t�QuQԛN��Dy��k��z{��1s~��%Yw����#SI(X�&���V����
��O�r��6h	-�����b>�~^!��4���A��;,�p��yme抮��#1	,*dݏ�{�6����v�y�ָ�l��ā�;o,�RU�D9ALD��k���i(�Ʊ����l���7�R�#5>�J��&��s�n�9#�ͤ�_#-|�"�踛�%~ �&�#�� H1�**M��M�WzA��v )%PrX�S�c>�j�NԼ�~�Z������Ͷ�l#s����ն���q�	K1 �w(�B�Ka��c�M1�{�&���U!@up〡�#���㻵�5V��窞nb�5�������dU0CS�)i�Y���7u_��á�ߧ�k�_�wj�w��G|�=Xᘞ�#��i�p�k�����^�뚡n��zbG����{b��i/t�d�O�`��A�-�]�9N�0ȡw��+{���d3W��g�J�S�gUC��m�Q�7]���s׵�\�Eb�8�xۈ��ԟQ!w��i�
����֒�I���piG�x|
�g6�����e�gi^��z�>[�A�/���aanq��XFh�(g���>��Kj�a�+��l~»6�BQ����!5�^��N����n{Bu�$������"�	�ZAlJ�����Q
��'�p��,$�l/h��VT@ص~��焌��������&H�U͢+�yaI69ف���>��r�,��_�#cŎK�^�7^�����1A��^Xs!�N��OR(�Y���[+Q�k��v��缂��\���N�8B�Q��z)��ĝ�߶����I<�ͧ����N"�Ƌ�;F粍E�}�q(�p��"�_�Pƒ�pZ���wT� �3�}Ё<��u���Z;Ed��00�`���ן�)�_k��:����j�ϝ�΃����z�S��4N��ߴ��B�� վ*��Ƿ�����b����:t�],�Y&��(ke��.`[Jq�A}�b���;Ǟ�V��/c�G�ܒ�E��[�G�ĝ�-lݠ >j+�Ř��,-�m�a�<����͢B���O1�!I��
W}9C̵X]�u�0��qǜ?�_tb�4������8�V
h���\��Lz<-'�=
��=I�lPIZ{@~Z*;g���m3{h�c�dt�Tr�p����)���M����S��xW`3�� �!��:lh�3�E�h�QN�>�N��A�k>���y�`4X�ɮ:=��S�������Em�t�-V���Y:��N�1D�'���� f5�;:�fq����3�5-Z�F�6i��(ݥ=%���å]�̝=��˚5��o���e�Lt�8�&�P��w��z�S�̀��B�3[qSSv�G��K[.�Hf�1��Ƽ�wgb��M���~���&@�d��L��a�ץS���ue	�����˜���cO���ƋE�р#Un�q����1���2�j�E��/)(Wz���!�?���3֕�=�|���kr�^O���f6�J�FC5uh��q5�m��"���!��Fa;F�Y���i�~�5d�<"�^�C��Hh�~E�R���X��;P�\>x���[%��I9/˕��W��Yׇ5Y��J5ɟS��j�N7�m<��@�3s��K��h4�We����y���>Z�/��d�Tփ#��nh�f(tw�$�I]R�Uw�xxL֩PX�$���k.�Jb*�P�^���v��߫!�ا�lgR�)��+x����8F/;蕺Mn��>�Ӷr��8K®�es	�e�=����P���5�o�̞Ki� s���u။}j�Q�Y�<a����^�Yvl*j�� q�R)�Է�eͽn�*����3��k �F�Z+�81ٿV����w�N��9�0s~��1�F��`,ҩUzS�^�*~� ���N���[X<� ������y�㦩�����V�� �(�nai�{;N>qIi��za��%r��o4�~�'��}�H�*�:�|�-s�T���͢�tI:J\�6��Wd���dC���(,�;�Wnn��W��^�O��ƃw)�	�I���Kh�BG�����P�=�k��;�#�SI��ݬ���e�y���Ɓ����W6}>�y$��%&�}���β��G�3+�RE��y7(��C�p��>���snM�{=�������mf��.n;��]1�����>g��{1>!;NF��L��=�bӸL�Dt�8��s�Tݠ:��	a`;�	�-dLu��A�i"��K�ةb<n1�C��dΉ��LRpfO��C��~��BK|�e-���MX�-�5������~�':�!O=#eLϦq��P}|��,6
�YbPD͈zc�)�&���N�I_�HΉ��#T�(F9�ּݣ�*'���6�+ۤoE�]����|ɑ��6���ǫ��:O"�a��G��g�Gj�$�ṳ���̯�>�r\U�z$bs�4H��C��~ P�8�`s��?�Ȑ4Wm��sQ��H�;[�kG�d
�FSʴ�G"���J���A�t�S��Wv�`�W�HXv(�}4O��~;X��>M�R��*Y�'��c س�{���D%O�.��l�.�/HA@��/��Y+���7�t�L���j����Z�V��<?���]�j
e
�A���׫	F�i�HJ_1��W�W�]�TJnI���d�u|��YM*�D�kX�W��v`��w�.(�*�����yA�CW9������	�&/}���R����֙��t^�f�ԝ5w�ʢ��q�][ZPr7�{���UYz.��
��`4�6G2��q9�H��q�20�f��/?��䑑���@������N�Z���vfò�ζ��a������ ��c=��S��J����'�EE��L�+�M*5ݹH)�q�e|W�Wc��B�=ܠ̓����6(0��sRTHԢ)��)��`:H_4}���*�L�+�Y�	��L)j�s�D����Q�@ �4fP�S���j�=��~�T�Ce^	�"7��a���,�r�(��ds*K>������tdb\�\8��R��p�����z���%7��a;�g������>�h+@�!��I/�.�ʰq�[�V�����B�y�ܡ������r��.������(u�z��^"O�n�3�FvS���e�^k�C"ೲ���lDFPT��W±�A��0=b�N�箹�C��p��t;zs�ߔx��8(��M�m3g N
����[��	H��5�87��'�)���q�M�Wc˅�hnr*<Y�F��cvMLfoWa�07!�<1�	�R�V:Ҍو�rb�(E�%<�ͷ�iP�oU��B��^H���+Ұf��vD��vp��uyD���F���b�gP���0�1��&� �ޜ�l�a��牲`Y�`b�H�� S��y�d�����p��/'��A7{�l�]KL$�ܡ�:���c��<|�ZF햛�@�n7&M�2W9��b�m<��͓�P>�Ptqꡌ�_����~���W >��mﲬ�����
��9��7�=#�y���~��ų��C�l�D�����݂&h[�S���ȧ���뗥��ɰZl���pm�D}�h�}�iP�B_�m�2�����)5����S��#1�YB�ې�I�]b0�����t�i�2�q7
�b��_0��ى��鞖�+���&����6�臁����N`����EY�|�V- ��>�����˸yr�gS�<G� ����3R	���">�$�����P����Z����*�+��(
�<a Ygs^�iY�	^19w��rf��4�P�s���U>�����s��7׿�
'�l{.�Y$:?&�����4z�� {�,���T�D�"��ҳ	i'����q�ګY�H�A<���!�"�ӌ�6���Z^��;�+F� *�L�u7�%�iHT����{L9����T<��!����2�Y ��#u�?Ŀ�:@.T �P�_�i�BԚ�W���/'Zqjb��H�9¤�&�y��e�-�9a�A�����0�2`	���[�b����p1�*�H�U����N Z�i]�/�j,ڢ4�ஂ1a��md�����QF:�%V��(7�N��u�ƖPi��4��4�J�ɱN���*�@�c���P��7�w� ���wF%$`k�5�9_���v�oR��ȸ?�oi�.��8M-��ǻ�ʙY7�"#sm�e0Q��hRnLp��v׽�.o��h0�J��?��C	P��BG�wK��$[��.T�,9�q��U��'V��~�^b%���3���8��c�P�G=���FL�'���8<��Y-�v��:��ݰ�j�u���=	o��r�[���CT4����"ĄAc�QF��Ї>�W�~0O#���{,��R۾Bk�+�5�q9�'+��a�U";�h�ύ�Fm`��8�QEX��ې��'�![���ǋ�*�
Х5Ф�U��z�z_G�-nׅg4fp���3������7���hi>���IFH�'w�7�<3����uΥ� D�(@�~泪�r�TD���}�<���3���p���Qh^"smk$F q����<�)��s>��.�Ɂ3JMQ��i�!:ݒo�z�xټ�A�Њ}ͳ�P�X<E��t�*�S�=�\8��).'�&>0���I�4������z�����܁Aq�=�Fgz�bU���9Eo9PB
w@�C���蛀'�7�.f��E���]7,jM�%=����ph�U�}g�2X12�E2�-̗��gæD�&{�1����Bk������=S�|����y�TE��w	>���11�0��g�M�{��"ėo^]�#_|C�B���/�`�h��Q�=�+�+P ��c{���o��>�T5PJ���kL����D��iD�������	s(������c��!��!�];]O;gwf�"��k��nA��j�N��w:۩��.�����"Ͷ�����5�]�w���n~�5-��\��i��Mԣڬ[R�>��%�=&g�s���YK�>�!��0on�Z��g�]l��=I�'���Å����Ð�<Ōɶ���	T��U���ZٜC��DB?~�<�3d���Y���;��ZH�U�ֶ1W~���#-��K�j�BX�=���hCÚՄ�"�V�W���8� ���v��Vx�;���#A%e�j� {�qՙo����Z���٢#"*i�Tz,R�b�w6{D8 �vKOk�p������	��]C��sh�#;O�����dP}��%��Spq?$�h�ɾ�gD�/H�)Ŵ�::>w��Eab��x���c��Ah��A���3b#B�3�����e1Vw ����tǊ��t"�6M'�:��N���R�Pa��tR�Y�-$��ζXQW�B
�	g��%��r���<"�Cб�ɣ���?h��[�EkT����v��o��'�N�0���a����u��7Ô/S�j���X��MO��	�b���7���!^��?��0��X����YX��wl56��^�sK�sG�T'�GT��Uh�%L)�6�WM�Jϡ�y�O���RӲx���m+/Bu7�������+��<Y�._8	�G=C̃#���r�j3pu�f�FV��8�t���:�*�?�����?�未��t�s� �J�ue�ykQz��O������D�_�`��k	橳MN+�FW�m"�w]-�|��8�Mc!u�`mB�STA�]��a��(!⮓�2n��a$��8����E˛�%�{��I��Xh\{�w�e6l!���AXc��ʆ*q����ƧU|	\�ZzT���c��0U�gWea�����!��O���/��~���G�ny.L�-�z��+��$G�L���{�ȝ{ǎw�x�`��_��U5�߻w�g[4�B3�r�����>���'���+E5�>���̢���x��4�M��oϾ>-�b|���tu����uQ5*� ��ݐ�.' %]�eV�EEfQ&�]�XV�qm#!MR�FU�p^�T�Tk�l�W�j�UkWg �て�Zd�{ܮMW����i�)~O�ސ�����������@;A�b��iw�h	:��K�5��k�۔`F�	؂�1�|�]�=y���x��6�F�
N��5�13A�A��s��G����w�Y���ǽu�E247����g� ��[�`\���'_��&E�
�͆��O��B٭��]u��S��[9QL�.��=���=���6�z2���>��^��dx�'�r���Q�����<����j|{����-˩�7-�&���v�1���Z>���#B�{������G|�� a��<x]�`�,)�l�o�������+��a�'��nEt�����6L����p�<\��:�sЋr����\���T+�����` W��oq|���������$8��L���7(�� �Ä��e��&��@K��p�����R���B�t���{��DQA��$���s����o
 ���PE�A��|A�������5�F��+j~.���
 �_O-�WI-UfO�ߎ+�[{c��	����F�*�g���[~iV�A'�b?ҍ����4eOR��u�+�lN�["CZ݀����5^�����ߍ4����n�)�T/�W3����.��*i�HӢ�4�4øE�򌍗	�A9sw�H�	��q4N�H��1�ɝ�~�׻�E��ƭ�z�fL�#���$w�T��Pv8�^C��v=�	��(W�� C�c�Aʰ�Y��(���-��p��#�k�tqǽ�ھDߍ�T�	���^1��7��J@|����~Gnp��&LA~:
=$d�)����GCw'r�7���>�b��;Ѵ�[{���o�v� ��T]DЌ7���_I��^@6׈�zBؠޕӀP�֦#0I&�1�֣1��~'hu&�{z�w�:�b	�����g�I ��h����$�js7# �WR\��٭��.RwCѾ��M�ه��Lv���H�9�&�]1/)�9-� �t˵ޭX��A����C����[#޴s�I@v:e�_0��鹻���������O�`wJ+�(�v�oBo��u>����K}v�<����.i�[Kɼv�xR.��)?1C�g[vϢJ;R������;�SPI&�h����p|�="Ⱦ�7���@Rj>�sr<h�WLC�ڳu�aK�[��<�+�*8�~e1m��X�M���#� Sy���_��Nh��ޣ'�l[���}m"�<�I�JP"�9��I-А�d��B�tzׄ9�h���R@bW)��`�
�����$�LuEB�E���ꀺG[ǾQ����.�̷r�Xq��j� *���+#(���+b�*��l��wu��$n2a���f �Η�W�_�F�5��vC��a
���Ǫ&�~a�&��`���>�e$ȿ���0�~���f
NV�̉�-gI:��&X�hߕƤZF�@;�f��F��2e4kp�����������|�WKa�!�E�֠�o��s���J�����F��@i&t�b����E|9�͓7�{T�i0is�-3AxO[�$�Rm����r_&uo&���EU�>�/e[{w��� |��|2��ğ��:|��#s�s������к)��a1��81�ry���<h��+��wW�L�݌��(3a| �WB���@��'�V�+l������l�8�>�ek?���ps���b>=q$�T�Q��Ɉ��Sp������<O*ܡ�IY��u��.�ml�W���؅�&@fW�ּ�4/���]�3� ��a�Q�2� �Kq�E�[8(l���*8-��{1K�������~�C��Mu�_��~9ݳ;w91V��0�j�ߕl�,�M��HEHT�M���*�c�$�D����b��J���%/�V-n��k��g_��I=��q�bo=̋��)I�^�c�Cy��W"2}6P����ž�X��Q*��GT7«Z��Rfz�~)�:Or�Qc��a�ױA��������R��S@rzJ� ��د8�Ə�O��˓�/�3�U^B'�7���Wh�����3�J��չ�. c��O)qq�?;$�����`%�	ꞁ�4f�Hxy��
%r��&`{���=��'RHQ�B�	@����5cլ��I��U�tc�{Y�7S�"m����(��Z@�iԞ|ޤ�<��m"N����*�l`�f���������z>��&&�ڮ����~Q%#��[��#�Ύ��^֯��$[��]v<�EBӤT�õ
�	��b�92H0T���)ڠ�AI�?nk��%0_Zqpɾ��b�l�*κ���ŬߐЊf��	s�!�%����x�Es\�2;@gW-G멅v��ߕp>w��K��F�؈y�]�������Bh���8�v�?(&��h��-R�kL��7R�ջ�`�hφ<(�U-h���0N���ȯ�����x�\��P�&R_0�� U���UVCÙ��$�7k5=�/O��lC�{6N.�pT  eI�Irj�N L�kh�J���l}�/UX!T0E�Iy�E̯���ghn�W�����a�J�ߜ��+��`�����n��	on��,0"Y&A�Xltq���X(�*�0~���k�a?<g��!<�8�UE�������ops�7��z�f�u��RnG�4�5�v��]����A|Ut����BC�s²*�%a]YP>�d�FfP����H�pڐH�YPqį���A��գ�3BA��R��KO��s?K���-�Y�K�n�t�¯@�!sz`�1�p�˨�A}���w�ژ���J��C�����r��/
ꜱ-!a��2�*�q����gX
�߉{�@��r���Qp4��EG��#�*%��h��"�NN����)���5�H ��؄*�d��9�h���!���eϏ@���p�x}��`:ҟhc/n�!�s�v?���U{H܇Po�����AU��鮙���(9���P=�;3gO}�~eӦ��d��/'p����Zk��2+6�H"���󎺀5�(?��zR^~��Y��z�<���^�\K@�L\?鲉��*Fv���&��!s�Kë%���Q�'��ƪ���ا�1Q��������Bn��[C3,!�)}�2>�'a�*���<4*��%��}����	��nfK���V�y!g6��&փ/�&�1�
�:�<@n�"���YãQ�������,BQ��G��@''���1^fS6�������eq���c�\� ��2p�&X��^~>c��Y��Y�����dU��1�|���ԏk�u�]�9��R���V�D�>���8�����j�:��dA�����QI�d�TU�|�L-�������s,��h�!��ݷ��GM�H�c|��f���5u������-	")�{�sSG%C7A{��(��n���}5��r�=] 1�B���9�1s1�kW7�f��]��������'8�ɝ���v��Sd��@��,]��ĲY���r%H�7S@���D}������rfPm7?H2�Ĭ)+�ظ����է��>Nڹ���n~�	�r}�b8-�7��> ����}ad�����vߓ�T�z��?���
�w���1ԤZ+�����Lៈ��/;��Y�T��Sv���7W"�q6��b�����F��C����v���Bnh��塦�9DT��AY�Eo�ٍ.�q�W���ť��`�hQH?��٩���Z��!D&�P��aV|�*S��ݳ�s�W&L��G�r[�D ��s��
p�u=)I�'7r
e��i;���Z_`�ԪϞ�-�]̗y��{a-����+;J�
�`�dƦi���=�?�> ��;��2������l��1�e������6�gCh���T��B��c$��T��b�;`3�;-A_��y�W�Ihؓޜ�b8;��QEb��c���KJO�h�Sv�<���:R�(}Ȳ�u"4�1���{>w��$%�b�,��xض�7߹>��n;>�n2 ���3�� �v[r>I�sҷ5S�PT\Om�a!'�1�s��H����P
"���b��'JY&S"��e5���>|��T'Q��bΗ����󎰷���욽r�����QW�z�lhS8d��ْ"n��t�e-Z��7	C���[R� ?���F֭h�-~�쩛EN��� ;Ƹ�\������H�Ln�B���o��"����\$!e���j��1�e��@�Dq�9FZ����w�W���1wE�w8.I#g�+��6��*㝽v�-�e�ߕ�X$�[��
z_۲�uF6D���<j� �4��0q�Ӂ~�NgA$3���9�S��C:V4i9?�(,�����Yac�j��GuR��LŬ���"��/�'�cK�M�sZ�T �Ӈ�9�v��ҩ��`� ���,c>�9ۨc�<*�L�	F�-��೰5���I�'۝���Z��O���M���I�.�A��e� ���.�#�<A�R!D�$!��nV;�u�X ��H���^�T:8OYc��.2a,��d^�Ӝ�q|1H�[>cX�fýxyi���',C	�\�ݓ?��N���\q��U'�w	�\��6C3��#6��ӹ��0������?��3�>��q#�9IŠ>/7�ܷbl� 3<7�a�j/Y��_����^�bw�S��1��ec�}�����H����,�CE��5�g�R���!��~�����
�Mt��>��rD����Ӟm��>�*�v�m.�e/Fq80NU���lz�)�~�y�٧�Z,���@�VΡe������z�h�Fԟ���c�/;��	y�vTZ��{��!h��:�X��|�Mf��<g'��۔XXG]{-בV"��?NgAZ�0Rn����9��@�J���i@Du�:|F�(��2(p��B���g���j��t��f�;��'�#��kOW?d��Y�,�����N��߽hhMj��������ɍE��Z�AP������w^��L�0���̌c��6*�N{��nl�/�>�+���
GZ��M���$�\���M+1�$[>e���'ܘ ���w��T��gZ��%O��;�;��?� t(��㠉��{� B�Iq��x�@�]��N��R?Ԑ^IG(������e�G��V�͠��֫tī� ?-HO�=;���c�[�H������;K�0���~āѼ�JX��jFμS���~�j@{���M�.�LBe�����=O����<�-�)7�)?&��a98j{�Kބvn�7)(]8�a6�A�9�|iV`�ʣx�A����Ǽ��8�fϤ#�2���,~̀���I�W%��h3�s�+�%�2�[�p�蹑���]�6��������ڷ�h��9���n��K�#�]��>jS���@z�"c<���+@W�����A��z����x�x���F{���?'ߓz�P�si����i*�,�	
��S -�e?���1�������U��wF��F�Ѥ_Ԅ�b�3�4��`��\�܌de�8��wQ�E���6A�h������v����^G�{F�_nMˀ �'�_���:x����6�*4ć��'u�_+P��t�K׳���x��,_x��0c��i�J]���cI��� �$��'�Z��� #04I�[=j�!�dJ��u6kQ��t��h��C @�Py����pd-�M6�V�2q�޿�ʛ�V�8�*��ho'�T��3}�ϳ�AдVh!�������E�6%��2��ä$Ό�R���cx.eMF���v=����6���s��w��":�"��\<K����č����gjL:y�ߥ����2kd1���܂&G��O�� ;����6�l_t��8G��C����O�F?�lɰ�|rs[��Lk7�N�k/���D-*k��
C�f�9M����	mO�t�2�f�c�?�h��HG��BI�ʒ�P��ߴ�2F."�W���2�0YȀT���[��(���P}����N�0��+N�"]8ZF�Z��ۥv�hh�������O���X>.�/͑c���;��*�{++nk#&QCZn�kHB�G3������~0���Ҡ3�c��D���0C@l!W�EE�:�ā�n�{A�����_���,���?�c���=��z	������hi���v8�9`l�_��w�c����c�)�Nts1.��Q2�ʴ��+��������[`A�;-)̑����P�tu3T��ꏖ]%�} ~�,.}P�(��0��������� �V$�q:o��4��zi�S���w�����-��sg�_q@QCi�}�-�Z���A #�Z���������p4 �2p�����&L�7G�,�q�R�^84��l!�Q!�d�J���\�l �;m�c}��l��(�,aº6�ZG��>�7T�\4����Ĳ�fŸ$�-�S�H�K-Aw֟M�6��B�I����V�^��ք�5���ω�N�-R@X��K�h�㽎3M�3��+��[����l̫w"W�C�3�����$��?O �$��oZ��pi�}�]��o{��=ad͝3Q�w�54��S8�9	0�9�Ҍ���%�c��!��^��X���R�Gz�`��7 dD�t(���waA��5>���{HW�%�9���ٺ��ޯ������K[��I?�,��z����0ν�r��I>��Tm��%.�9��1PI��Lu�1��s�}5^>I�7��G�Mԗ9��Χ'@fX��0�,ֶ�����9�%�,�M���)4D�h?/ ��b�]��a�|'�?x'�qJ�"_v�= �L�H�q��k���x��T|()�Zb�sH�ʂ��r|�n�WbZ��U��M�.A7�w;��V9��6vuމS.�ӌ�_U��9a�b���|omW:6G�@�S�NB�˫v9�&� 5=��4q0�iI�#&d�~�j"�"�fE�NcR:�vM[����8��ng]���B����\\��s*��>�݂�Sq^�<9�VI#�\�I��upU$�b6q�v4i^�F�;�4�|��W&�u���h����S�7hk���_�C$�C��).%�͘��[��R���wһ�r`�]����l�&�s#�x��;r�<�VS2t��]��5Q��|xF�%��a'~|~����e�"_���5z�eh<� ܺh\�;�+~#���ϗB㲁3����k:�TZ)Ei%Q|Ac�2��fS���"	��_� ����K�g���h\�r���u��Qq�rq�j�4�!��ù�S���w=;��,L�cuC��gʕ>�y��oG��(;���f��;�l����u�y�IK+/�8�KKK�Ѧbi����NcI4�T?������+� ��F��D�x����w�2�lֳuP��_�?�g��FY-d��2� ̞��`�Ѕ�;/5������<B���������SX6kN���4�����;�2�d(��NoU7���#Jyk�D��,�Q�%ߨ���ߕ 7@����xw�j-�o6�8?�'I/L��D[�*$lY��a�Y7
�y�6�j[��{��k�Ts%2�B�e�3�$��m��M�v�G�R��1�#5��N��<=��l�%�	�N?��^��'�5�$T%�*��N���W�]]ԩ�F?x,8'�h9u��:�=I���`9ם�o��S��~��r'���Ӟ�8O��J���W��<ȏ��>$a[>�&�o����}#<�\!�6���]R����]�{?N�b�� ����2<��c��o�\"�����ĸ|DqnT��x2s���\�d4��1"@��=�~g�E��z{kGFy��bSȦ��L�����a[�����72X\����~�R�B�ԧ)��y-5�W{CJ�3�nȇ�����`�R�4�\�EV"���_�f0R��K��+J�F ` �/Ԋ�ik�ݽ��pQ��5��9Uj��
�����~t�8&���!H�Y���6F��e"���` Yo��ב�a�����'��
�I�`�)�d9;Ş�z�I����ⷞ�d�2|�CM�7&7?�E�v��9�y
3�p��?�C�BP
����s�6�m����r�̛vJ�D��p!����.���Pq�1�{����$���l�#Mn�*ipkp��уy ����� ��5���0�4�Հ�y���]_6`��_-5��ф�5(D͢P �Y#�勚3/����:璬��)��ކy����ݒ����-���L@Gq��`P���?"��ū���Ԣ����$����\�݉�A�|���t�!��>Xoqd��Q�#ls��{AZ=�޹��_���7�����9)�Z�c�&�k��ػt����v�"0wG�G��8[��z/����K�(('��$(�k�\k��C�w�����7L��S\��d������1�>7��~�d���	
m���j+�mȐ3�<�����̍7�b��������p��)�X{�o���@�j�-MC ��Pc��o�BSb}�䁫��5�F<V��%;�ݳ,�؆��D�����a��>�ƭ�l����.�)E�le��Bf�YUv�BX����`g��gˠ�G���:��$�D�-e��Ȑ��6'��sX��f?���,��v��Ob(��{M���ߊt�*����S6����iFnh�sG�[P�ҡi��MnH��O�$%M�:)og�h�5V���O������ܿD���q+� S;�1A�?�oՠt:8v36x�`GB\:!>l�e�P��Gn������f�&w	w~��]�{��{D���Y���p1ϧ0�����c][����~��A&
���:g˗��K}�ǅS5�+�69��O��}e~=MX�0�֮<�R�b"V��j�f3u�Q������u��y�i t�	m7��ݾ�:���Ku�i�$����Ku�Pĺ$�|�������6w֝��Ƒ�8hVܼ� t�w<g���N���#�Rk�V�~�!uo�]bF	���%������wS��{���T����Ap?N���#� U01�gb|��N?�5D��.��;N݋א�}�y�$_D�FcW��"���tBc*$TtxPz��ʄ_�&(��GK �%�272�3I�����$c�Y�sHm����E��}�.��2*�*��[�NB�)"U3-���i	g�n�ׅ\�;�q7�$��Nt�f'��b���a���R���z_�����J���`R���I��N�N��� �vL;53� �nN˸/�8,1����ҚZK����)'q���أ�h��y��.�5`����"in��՘B:�����8���4�x�zzO�U���U�0��9��E���`"�+��1��*��������\�Z@�%�P�����F��H��z.h��҉�R"�z&�.���z�m�g����;���c8(�?v!S.�HKde,Q�q�wJ*��X�����]�V�Lv��ZE%Ƞ%
\�����n��T^/S�{�-{�����W��B��c XΐX�-̍�aĲ��T2�g4�.k����d�N���:��!���������!�r�&X����Y��8��}I�m�=
h������b�佳�����
�^�PW�3�mI�.��G{��M�,B9�f`���q�Ĵ���3GCD��Um"_�@�Τ'��%HO��ğS�FS���f���jA��F�%�	�Ѫ��@�ߞ�9�����ԉ�Π=�c'B���\%ڌk���R�Zz��)�&"��6�
�_��,�W��pZ��q�5�=�Z��;�&�'k0��]�j���S�̴,�������������,p���v��hc]:��[�F���.�$�z�O�D�"Ecx�˾C(���\�)Yr��+2����K8m�{y}Q��xis��n�UI�����-Ұ/>�(�c\��ο.1��z��9lї�z�Jk��լ�t��#:U��	��[�+��a�<v	G5��c��e����zĶ���"C�G�1��6�:���1��2��A}�M�z�i��Ƌ�s�*�Ū9�he����L�̄���S�������^k:���B�PJU����}-H�>���}~���xf�p���������<q:
��V����ո��_�����$�#c��<����K������񮑪��}]G!̢�9Q�0 Htt�2d`T�>`���[r�y��N!�����7���vO�M��/t�;ɺi�s!�]-����!FU&zH�m@����Mo�E삗�"��R���1�"P�W��=y�����5�QqJTa���<'��L����4{X�͓(i'�G��1-�3B��v�~��lha���=*>:�$�٢k̻��#�Q����=��޶N$%=��{=�{��簜���b�Y=J�B���qc��n^�cU�N,�E�*	 �w���%�����R����ȁ���@:�S�a%-l6�F n]�xr�)�+�)bו���]�3d�u@���p���������
h��G"�t9ĩB�^�ժy�+�#2��/,}	sY)�4���&�Ưz6�GRg�rS�ܽ+<���&�X��M���[ƍ#V>�B�t�7E�󤦍�qlɳ3�l��cF��1ȒP�c�~ܱ�"�F��9�b�?�����#�l��};��p�q2��i�ϴTԒ�+�e��l_�w�)Ⱦ��I�b�i٨0�ُ|�z�g�c�ϲ��K�it��.���< ��Kn�f�/�Z8���.�����w*�:M��>��ЙnS�=�=�ku�6�S��ea��\b%x�.l�@�Q�D��T��_^F��� `�dQ]����&�D�@��;Ag���$���ͭ7�s^��f���8Pɮ�T<FޑU�
���3p�%�w5�r�a$3Dj�GQ;̼�KV��Iq��z��
��d&=��0��o�Z
�Vz���i�[��b*�y�P�::N�[(!�Zu�����d�=eo���}Uv�Ӡ�	�x��bU=���ޞ"����!�#��ԈQ�pC�tmFIR=ߊr�t#�|z5�G��Q��PM�[�mb�F�$��:��-��V�ӹ�,����/ܹ�z���e`�F�}ƴ�B2�nF��YHtٍ{���2 |�/�#����j�s�
�W�_�@3���2��@t���tR�	P`�Ρ.�l�o_���ӟ�i�њ����d�����; �J�L����a�d��YADfdl��,��'����h�	hn0�e���2?�>�f��:m�
�c��I-�:U�&��0HX-�����h���k.}�Ij���oo����w	��WD��˿Jx��75X:�"8�W����ԎI]~1��T�5c�d���z�����p�JR�o�M�z�".��r7w�W���$� �R׍��d���^�A�����do�]�"�nf�f��ޅ�H��T�j�-�sFͦ�2��Q-�����]bB����S�^���&�d�=0󑣏1�5�^'[�>"�P�L�6�F�; 邹��T�^W��G� f�M�J�>�Jot��Z��H��C>1���f�bT���\�� �V�jV<;�Sd��o����NR?��sb���V�>����^)�"i���?3��PQ�w�1��*��\�c�];�-���Z5��&1N݈r�l"�v�+X�Y�\���/��c�9ɽ�梙�������P���朞-�wR�V�e}� ��h8�,��h[&�,��G҉֠[ޮ�������e�[�����~j��nqR�S K�����ElG�3c��_8l�G�[�9�e�:��oGv�,)���G��R���E��j��Q.<�?����(\qh�V�-�Ƭ�3�<�L� ?��ǎ�x&4ٷHF�w��o;�ȳ{~�����p+����5��N�{<��k�3���e��H��x|��B�_�w(�m�����b�������z<D�����W_��zr@W᫵S�W�����{L�/H�8=���2�h6�A�2[�1��l���lPH����O�]U�#§sY��x*e�S��<����v�,��||���B� 4
^����qEF��V}�\{�Ev��]�-���j'��%k����_��꓉��d�K<0��f	ʿ�d���l�׺��� ً!�3��LmX�h�s��<j�u~����t�ͳ&�7q���WE����ܙ�;?�z-�^_�=�!%����4�v�;������n�ܴD�7(�Fc7��Lp8l,;��D��iJ��|�<��Z�8j(�e�	�FwK7��׾���c�u��Ӯ-�
�ōp��D�$u2��S)�T�������efF���	�Ғ2�1SB=�ͻ��)O�?�
t���u����Z�,P�[N�yW�d�t�"�R1�{ �˰t��[��d�U��6��9�[Mx$�b�ֲ/:��:kG��NJ��úXև��Q9W˻�h���$|[a��A�v��1�B~��I�����e�k�N��E�<#��{/�*��1o}RC���l`�Z��md�D�RS���4H31�Y�=�3o�'>@�x�b�Ev��K��� �˃!�?�q^�Al�5���2����V|zѸ�rpO`K���R:�vh?�HvџXo�e�ԟ�=]N��w�>vh/��
����Xwl����	���4�I̼m���T�� ��(:c��1�D�{�J�J]�T9N���^��dY�E�T�{0}����v���v����|I��9v�XDR���*�F�J�n���Hu�W�z���81�2y����E�a�K����˺C�����:������!�~�����L:P���R�O9���2~� �'��	�<���
k ,�m�oN���<0��4��@�/��lF�&kl��k���b���\��ُ��Ji	+(F��&o��ڶZ,7,~OE���o�+f^�n3��7��[o/WN�̡'(;��eŀ���&3��)i��m��>�t����9pl(�&�{�:�1eyI\���2�4�yDn$}��#	���D%������(��l������[����-K�����\i�����{1�z�>�r\���g���
�=��mU�_π�<�1�������
c��֊�X��U�>A�+�.>y������oCX�`��k�62�a!r��kf����.�zx�L�I)��>�[����o7��~L����IGb����S�8�i�n��l�P�{�&��lK��:9jjD��/��g���a�3>yk�"i��%=x G]>h.��ܯU�r�ޓZ�Jq�g�sр�V@�Y�LeB�����ȱ����5$RKè�d9V���{uĴ��l��2�U�#��a��k�6��0���E�$��VRt`���m}��D��媲��m��9?��{x�I�^":W���L�ǌ=���<T���4Kǖ�i�j+��Ԥ��T�{�g�R�ծɥj�+k3��ҥ+�z�1CV���nv����;'`�?�p�-+��/j�_nPfo^XV�R��`��a�q�\i�y�~s,�l��a���~���Ñ���ے�E�T�[^Rp�C�j�3��PP�QW��ة����9t	����u��>Q�N^�͗�y�߭�=b�!����パ} ���v�ɠ��9���HN�Sw�.&1�f�dSGz�㜾��*)��F��^�OP��Z��(�:4�F���Hj���V���%��2|������ʸ�`?Q	��Dr���,�M~2��A	�����Xi�0�|��q*A��'��d��Q��o�h*I�T�x7->�(��"�G�=��%~|,�꧀���yͷ%�����l\)��Q������H˩w����y��$Z��'�G�hTp��db�7sW����/b���g1b��ױ�>pK������[(�B'�F�u�7� �H�]�bZ还��g�/@0��o����/�q�n2�y���8R:�([�c� W�}(4�����n��J�6,�7�!��X�����x�؁�K%�;����s��F'� �6i!l�\�_����f�`�ԽQ�(���cQm.��b�]މMY&8;�=���9l�p�����h�=HIx����^������]Rj�R���;�W���G[��.���śK.Ę;}��[	s�L��v��m^���{��(����,cLU�y
�֖�����S/`0��AqC*��0�w ��08�����>���s"ۅ���퇑�7�e��H���%�
&������]޿I8~1td���\�fZۃ-w�:�ƞ��!�����գPkww�Qّ�3�ИF��t�q��T�᎖�;�(.R�@'�MSV)Љue���=���d�P��A�K��aka�\|��^�B' �	���Z��d���7F���>���b�w�?���K�QN1��'�l<=�z��S��`���n���8@�ږ
ʽy�Y9�c3���"_��Q�vp&�����k�&ah~cab�%�]w��ޮ�A�;���v�"��Ͽ0�FS���?�ۢ�Z��!f1���gv�����O��XѡGt��v{b m�Q�/\�e�b�j�8��M$�&�r���4�4���:X���h���{(]�p�ZE�:X�p9)Y�q.�ں���`)�� � ׳P��nE�g��/=`�U��]&wJv<�U'S<�oG|,��f�~Tw�GR�\�Ha��C~��mz�i�m������ū����ڑ�'�_����5C�N8��=�U��F�SC�4�g>�E9�!�&C)�H� ���� �x��PA-}^�:�A8�z6�Bw�{� ��<9�𩰔M� ���Φ��.������ڒ�jH������q>>���ئ��U?���~�87 �m��X���`U��6$������$�F��p/����|���y��niZ�E�,oPv���><��)��،F�L���EG��a1a]P$�L �&i�ZK�P��z÷���5��{(h	���ҺV\Sތ�)C�$N�,�\k:���b�D����ɱ���"��J�8e	���
���20@٫�K�dx^GǕ�R���9���F��k^�qo�Y����s6��yO�
~}u(��@��άo�v�q�q�+�.�Z�������<l�m㮝���a<\�V�o$�شE���
�)�P} �������MdtSe�p��`L�
m�'�,�Q�\b��X�zF�4�T�y�!@�D��F�S�V\������KU���\��
lF�"ߔ}K��;GE����紞��,��=��t���E$�%Hd�5�Wm�D��u�@
�A
r��.��RK�Q�cB���������!+��R�:�Lԫ/~;���Ar�3�����	@͈�J�?)���ν�>�~|�ݪPs׷+�\r#�G�S. ����x����(q����/�
B��j�ذ�3ޢQ�ܶn�B�DC��	��ϊ�Zj��� 3�H*&�<�:�q�U���:���R��m;��Ʒ0bcQ���X$��a��Som�j������.9����+���:?��C3�8j�t� �3Z�m �N��/1�]���d��6�8�&�y.(�s�H"�@�)�n�~PL,���[�ْ�|���rl+����$S���\����Cf�!�YM����H�ð=��E�ķ�(韲���Ye�����62�O�Fǌ+�'��$�nʎ6Yݒ��Y�8����������e�gi��F!б�;?���0*G �iZ<1K)��^������)��`t7��Y�h�~�M!a��]�o��߈�֫wɯ7���͢ICd\����4\��Գ��c������3p=e���\`r]�y��5��E�6���'�W�����O���Ϛ��W\�?��@<,�nWzT�W4�'�ȳ�t�F��Ea���G�-�-AN�5�$&�˧�9�o�ê�;"vQ��0I�4�8�:�0c��9�����O�uޡ<�B�����`Q�8>[i�_��p�"���po�X������ӫ�E�8�;��.�돉� ��-2J��T{;�n �'>V���4��&+`�v�GF'���σZd�?��>��;H	�pv�4��'Nd+ZX;6�wh��J�b}�����|��$ZN�� Ћ�2��K�R�F�~���逑���z�?->�įL����i�>�H�7�DhPv�j]w����*���ϖk2=
\s�Z@�UW�iN\UC:9����_�K��	2P�X��b�	o>��[�4X�au�����ut�$��qĉ$�f`��7���̠ ��ކ���Bz�X�y�Ѩ�95?��\,�\�����6�T�[���t>�V�6���i0䙗��`$����d=^�`��FNZ1'\b{86��n�Z��ns�Ц�n�I���cXO֑�zPFѳ�B�E��.jJ*����<��"�Zq¥n=k�7.[����4[����`����S�GԂ�b	�
>�$����B�����}�Ȗ)W�y��N�Qٳ�����ta�R���[�+�]�r��yk7(F�|�֡�(�R1&��7`�1��GT����S���iq��`�KE���i����r,�J���=�����R��I}�ŧ}����[B�LZ��ñJ�s�U�w+x��M<1����ֻ��Czs�e���`4*�G!�����l5u��'YC�b��Anzv��kC��7��Q���Y65���s
6Z����GFa��j�sg#sՎܜ,hq5��r[^(�Ǉ���sP�v���!�N���Lvh�J�!�$�#��y�a�PyQJ�j��L�	�\mˑ�}{q�6���:Ǩ��Zm�.���Fo~�i��0�<q��m�%u*�S�)��J��D���1V��l�Ѵ�t��Xpŏ�H2<d�w��FO�-Q_!Jޮ��QX�<i.X�(��Ta
���a�)�~6�f�=��]�MH/.#���
���E)wl�[t1����Fh������dD�)At�;bɳ��k�M������"T�R�j7w�uq���⒄���|��]�}�{S"<8T b �:����T�	T�l�����yʡV��F�fi8���f�j䳪�Qr��������A~��\]:S�g��]*@k���o!֡vҎ�%������Oc_!��H���%"��:�AwN1DB��;��S��S�[�-	�+2�ΊF��̰F��Ŧ���N(E�~Saz��`�x@3�j���MF	\5P*��󹐏uF�_g<��R���͓�,,IC�~a�%�IV�=�j��n���-r�}�,�����-Oʳ&�'k>6-����!��iY"�xY�<���.1?���#��3h��9�a.X�8��@+:r�^����)�"|v��si�m	�K���أ��M�W�|"�0��u��T�=�YN��Gx=,�G�UkD[:��	�&*�ń��Vɸ1�lQe�)޸:�L_b0,�Iy^�y�����?Qx�����b!mt��)#Eۘ��ʉ�Ү��->(^���\l�'*(_�Rz���몝3Y�����%1���+&M���~�ݿ"J��O�΁"W���CK�P�K	�����6��킻,H|t_�"���8�#��J�(���ν
V�?e<�;I�B�NRA�
���s�/�����s[Z�E0�����-��zg�,_kx��s��A�pcS�k댕��u,������:�o���@��%r;RN��*-_rpX�_��rؼ�k�]V��Qx!P������"�=��%��+�?���(��g�'E��v3���	�a!�t<�w%'��Č�KwE�Z�-���t�_p��N�;^8��ߗ���A��-y������gX|�$�{��/"���ީ�%�����͞Z.>��ϳ�PY��]w`�m����t^�^�Ƞm���x(X�*i<p��2�2�_9�~I�)���<oypt�3���� ��ʶ�ʡ��������D@#c�����NKP5���室��R��E���h�o���)�f�)�3+��s[%��	+���'����E���=HfٜD��ؖ�f٧�e��oG���J�l䃪�B��ۖT�	��6^ir�Y�90����	aiV�:�2%��R���Z��޿��h7��x��̌1�E�V�[�8v�}��T����Ѝ�{C��=�� �V�ظ�Am�U�ה'6�	u��:��$9��v�G)�E���k�g���7m�v�
�+ 櫛���Pʠg��@�:%�*��R���7�������i����jʪg��� -�����"˓����tX�"�V�!Ѯ�!�s+M��4���l��B W����g@f���N��-6s ��5jiU�B'@��#d�J�ȵ�֢l�����7s!������2�ï�� #���^�Ϊw�0 ����;]��)L�g;^C�;�-�e�L��հ�q�ט����IU���ެ��J*�c�$3�$<zD�(��tT9N�<�Jr2m^����(l<�4�v�_Z:i����Ex@�����m�������E�)᤮�ƌP���d�[dK�KTpZu_{�-$v���&:C�A�rо�J��t�b�r��ZtԗJ& E�f����m[���_���w�s�� q>�������v��2��p<��I���+*�4?�H���>�{GA��W ���o����4u%U.P�)1V����_{�6O*T��z6��i&�*�U�j��wZ5��]�J>A�௵a�r{W!�2�c/葎���s�X��B���	���2!�&>ﻠ܎�������AE���J��oSs�q9=�5�^\�·���mh�|�ګ�Y�i�_Qja�Kˡ���Vcn�f���i�M�@+�����+FB��[�����K�,y�:��� ��_M"¾چJ��u
;`��a�F����=��:�� 9��5Y�K����n6��5������̗'���<H5�n��ty�)�� %.Di3=�U��)vO�eA��-����1��<h����5[�{�4���J����q`0�Z�dʅs�Ta�2�X=Q��\bS8%}�T�~O����nh�Q�yO�9��8��YV���,�5��Y02�
�t
5�����nMh�J�$��Z�`hZW�n�Vk���]ޔ8A��w|�Od���>������׮u�`#Y6����B������IԄ2RX��i����5�:m��E��Z����qsu��zt�Z��Q�m�|����K:X��@0��E:��u6z� ���u�����z�#<q�����%�q���,r��C����.���ˁ0s9�����Kk"۲ס�+�5����e�r��D�r�q���XR�(�Mց�Bj���!���Kd>p̶�=�A���۟�⪀�$L-�{!��@nƐSt��Y].Z��.�
R;��$������<�����獯�[��qb�F�A�?z���z�N^+���|����T(�)�3]�6)$*! R'L�x��D���w���ڇ(�&��H���ʹ)Vk����͚�/*�S�D�NA��KH��m���ǡ#su�Ӥ���������͕<Ehy̔e#5z��Z�N���ܗ��4VY���-��S���8��I�n��,�������AX3O�S�(T��dj����R��Z��8�\�$��EW�ŽS��G��wnn��:��i�F�\���LVW����1���X&�m���i�~�Z1��9S� 	�Ŧ��~�ٟ�(�#<m��^� z���s�+TI�	{�����1Kq�_b`���F���!��S��TR>xe+��)]���*�s'(��}3���x^�O�����.Œ��`9�)�M�ѩ��v�l�u
x鞱�ڥp�|�zAy�Wpa���0o���4u�m�F����<�<"�g�E��A�9�8��z�n������@ceEV�DڼS�[4��y��օ���}�o��r�8AuJ�	�{hBs�>��*�n�U�`YwL��hK�D���`�M�Kd�b�͖Q��R���K�]�����>��q-�jp�VA��|Qڂn0w�m�ʷ���
��Z�BW�ݼ���{f)�(�w�]�&|�6������Nm��Y���#�%f��i��I�[�a�v)��L'+r�0P��ƨ��Q����=[��À�0ӌ���h��x�e�F���W9�M3������<\�-���k�F�)���
3��%�Tf+�3d�Ԓq���j�����Fe�� o����h7��h��+YҊ��T,�Ïh.�����-x�<{m�c��!�o�����XN���L�"�6Y��}4�9p��]��Q�2U�n�RR���?	��;hˉ�1��Ե�x>&F���Js҆�.	��;:���m���g�5��,CZ��5��C`a�-�.�Gvf�x�3tf�$$
P�ʂ�c A�إTsx�s��e�Zɽ������I)����nU�����5���/V����@�߮�@�ǸohwU%U/e�lĸ�gP��xxG�$*{r�+������ ��
��,F��9\������A�Ư���J�Z�I�N��ζ���Wː�C9��Y�~ ���z��r�]>�dȍ!�٦�2�^N���(:(����Α����qs�:�e�\�0G��rp���VF�<%�)�AX9�<cT^���b�r�3�P[H��Q�u�	H^����$Qu �SG1��5%�=k*,� ʥ���:�-m�����w<�k�_��<��^��pSj�YV0ɘ z��ڭ��Gd/�3"LU��Q�ƬΧ[nT�9U_�&a���K��ï[+<{���`)}�=��$�I�Tˌ�lR�_�˞���Z�b)nk��`9�BBN�m�f�X8z�j������"�}��ݱg��En;.TE��vjm���>�� �x=Sӡ�.c@���䡱��xTՑ��g�˄�6ΙT|�t����+ֹƯ9p��α���e�TB.�#��mnhzP%�pbc��^e�|��m.'⑼��Y�=j�!uw�W2Z�%�,E�����|�^~��f�,�M�N��i�Y�����FS'��h����F�]�L���X��������TUR���]6���4
�k��򓣚%��\�@,$`���N�y�t�^�<��2� O��ދ(l+ݩh�h4�Z��2{!�/D�f\��N�0�h[+g���;T����Z{���D+~̕X�}qF�5'�����L�ݮNѶ�XO#M^*����L�.����mr�9���J$q�֟�.���E�[g��;����+
��_Q�G	M5b�v��g��.Geõ����.w<�_jᅩ��ީ�#������n:QJ�Kw����ȓ>�P�xً"y�uj)�6qъ��u�ʦ��=��h�<^�(�e���;j~;-P��z�� R�*�Bw^Q�?d.6�ｔ(�~8���6� ���w�V��:۸-UN��H�ծ�L�~��(]���2��<!����ޠ��:̘���h���k�>;�Q�4���`��(�(OmDP�����m�?�@ͬ�����>E8P�pIA���&�� �i��hZ`ޒJ�ĵܧ������qv�|����ᤦ�W�G�sw���.Ձ������t�e�R`�dM�+�\a�J꿏��6��$28�����1`yg����>�S�� #��J�ӏ���:OP^���+Ҁ�ڙ����l�m#��1e=·u�G�h�`v�$�����#x6����mm&�r+:�k!y�70��irF��w�m$��hNFd�w#���(�|�|W�]���3�8	M�}����q��r�r�Fs3�X�C��փ�TA�_ArX	���xp�Ғ$�G���P~it��)/��uB���g����┈Ĕ@��֋mm Q0�C�s#)�r�#��'�iWs��t�n��9��"0��`�dD�ѿ����l.\V@�5��'�kJW��!!U�ʾ��3��^ߩ!�x�`�?؛v�w�_Z�G��g���;�m�(+J��q��X%��E�t�'��;㶰��B�؊�d��/�"�7��Y�!//@A����L�)���z�j??\\���Ǹ�%�z^ޓ\��>�[���2Q��z?���L��ȑ��"�J���ݻ���A�� ��.�_s�4�C��j
�XA���y�H̦��η�"|�������b)��s�XY���)�Y������g2����Ǭ�͌�z���|��ވt�ZȻ-�[��v���." H0/�0��	��Z'2��c� #J�%a����M�G���
 �U���t�=a/�K.}}�\�%�s��a�0{Kƌ�{����^c��2W�F�t��_���B����z�aQs69���4���]�}��8vp�(�����O����L��-��<������� ��4`xYy͒�T"����%�u�&�`���`�14�>�b�my�68�HTx֧ui�J���Vt隨��>�
Y��"�����-��#�3H�M�Zb�E�<M�J��D�n*����G�����5k��:�n��|�ɱ3�{m�R�C�4,%�!�U�?v�'�?������^7u��G��kG�/��mY�xG<RRzY��˗8٦�g�U{���6�6{0I��U�+�*Xds�ў���/\d�q�d�w�V�����]Ғ?�,��9^�����a.�8g/.�F_�~�����M�A�2`g0��S�� ����H�X1�r��l����ԱZ^�Lu�]��.��W#�8��'ǈ���r�����6��?M�bRψ�+U��7�g]t��c-���J��AS����%�?Ϝ!ߧP�!o�d���R	ʝG4�:��t��Ao�e(����Ѿ�iS��������������pj�������ĉ��L/�K!���$�v.q���>��1��Y�z���B|�^0�������;�Y�X/��&$�5ԗ1��U�4�����_D2��|=���y:��S���hy�Ka�h��DW��h�6����D\�h�4�\��b��8�0"�{�(�V�@H����6mHP��-���O�Z�=�@k��F���X��$,b\SQľ���}f�w65�>�:!;}�.?|���t
!l�Mن���=��d��@������KtMFmӀ_P��Ndj\���>6��x	*��'y��S���'����A���w���YN6�$�o+��+���T+��9c�<�@��_e�OK)������kK}��r�/�;:�2[�å*4Ӻ�j��� �����
i~Xl),k~�-a��	��_!mj{�I�a��AC��ŉ��kp�AO�M�s�:�~E�%��ݼZ\%O*�Yh�I�6E/I��IY�����|���%i&���y�)�Ҟh̥E�E֩[�4��-#��	b�v��@\�k�T��� Q8��*4.��p�q��[��B��7M%�#QW�]�4!��$�C��ʍu��Z��h�(��F�K��y��[BZ��W�c��%�I��{Q���Y��C�{D5�C��jt�� +>d�/�{���CR��~b]H�(ٗ�	���щ��V��ր�Oj��4!�+���
`s��y���H����F㓽Ӓ��8I%��q����������)=�K�W�sl�
2��Fݘv�{�
�x�o�Г�oо<d��+�g�ײ���Z��X-g�@�MZ��xd!�������'Rvǰ����|�fR�� _�Ё����D��s+m��e�T��E���?��EǨ=����M�lL��t�uW#j���:w�S�Bc�'��~�:��Z�i
�C�9�s�jG�ޖ,�=�yK����ܫ[���m��y�KK�t�!7=�3��Q���vvL��>�d��%Vè|
��Q�'�Y�m��^��_����~W��l�#E�v��#[�z��3���TW^Pw�N(TȤhc{�2�d�n�o`꼲N�p}C�74n������x�ϑ.�H��Ѯ��'T�9�9?��0�C��lJ�H�xl��v��#f۝@�|���&A�gQ}i������#A���+|⥙J����.�O��V��x�9�8�2#d�͚�0.��Е<�{N]��������(Y��!�!��NB��6 ��"�ˁD<^5i)Q_0�|v_�s-�rm'9P�R�N����}
�Rw}
|�� �Ѵ�����i2Q$����h�G���AC� ���3�/i�;�*��9"eS%��D����u�]���O�;��<d�U��\B
e^�sM�o�� ܚēB��%{��H��1�)����H�G��j�cD��Rra�RL���N�ёA�}�j�;�,D��f|2�W���N���%��K^�+�u|�&��'�I=��&��q|� ��{�?�����\���8d���|����_�s�f�.���)[(t��/�ly���vO �TU�wz0B�f/f#D^F�,{ ��8��X{
m̑�:�u��	#gm�7���{B8]ȃW=��Kl�tl���(L:�U�=~r��KΦ&жHcΙ���)+���Պ��6,��w�*Iy'�g���?r}Rd�FN��`�������y�LgZ��"�D�7.	y�j��)Q�M|vؤ�މE��ӥV�m��;��ǻ��#C��4��7C�B(A���2�i�6r��l���c�� =<���/��c��c��
4lu��!�
�y'����~ݛ��F�F|�n4��
t��IZd++��H�L�D,U:��w������~_���!PF�J�=�ӷ(�|��'�-ǹa:�����^� �y6�>�-I��ч��f���xvh�[���&�*rT4�(���w$����^s&Jր'���}F�W���Lyv������)�Z���Z��A�k��f��T|��g�4]��(<j�}0��Ъ}QRK�@��1#�N_���9B9�dg�O��]�s6�W��f��f�d�O�����f�
[��]���m�) �%���3�X�����7;��+��.��]����yT3��"�ob�h��}�;i.⯷�?~��C��-H���.��ݬ��Ȭn:�?v����b�n8�%�幇HT���?n4�$���X0�xK�b�p�O��Z� �ܔN�R�&I/�K5�BM�tWD�M&Ǧ��
����SLS&eJ�:�l#A !�G��970*%�fr4�ڗ�2��ȟi���I[h�)/pT?d�<(�5Ɨ:g���i*��*8ڵL�Zn�:�めU��"6��V[��
y�Tm58|�e5lT��FO��Ƣ���{n@*�ܖ��1�����{Ba�Oqס
��Ĕ9���v������-�9�d��<�G̎?�r����af����	����#28c#S������Mi�1���0>w�TeL���(Z��Α�9!ŉ{�������F��
E��T�4Hɧ+�%��B�I�^���}���6"xL�
NS�w!H��D�-�*At�=u���� �Q+�rK0���	,��G?tU���ȯ��	8pq���8����{��z��G:��;�3����9y��sg�\�U���9 ��p�#���Q��I?�Z򟥳���1^8�}�r�](]@�m�]��3B���(��؊h�?a,�뇭F�����|��z�6���tv����|�^�b:ĝ�Be�ei�33�P*���Fky�c�F�,�rh�7AZ�c�yL'T�٠r�gl����2r�k2 D�?c��9��s�WPA����o���ٲ�AAm��=8c���r���2��ÉQGW��|LI]A�̃+����I'עy��g�=׆9����4��7�i~�Ԭ�j�_��$)��X��ˬ��b��I[Ô%���̥~��E:�i��
X��zB�O3�nŔQqb�Q���Ƈ�������ߋ��waƄ��H+��ފ��(��d�.R����n�hY�S�k�6k�	�T�*�pD>%8��y�V}���W���x�F:����*���Wcb|��&��*2�0���8 �>�
k�vkT�mΉC4-'�B���?˟��~H��Dn��i?����Q��%;-]0^�'@6�j�?�h�^���#��w�I�q���8�`}��1X��3��������#��hO�A-7�R�����agwb��ʋ�o�G�!e��]%G�s�*&���+Xh�	+l?��9��f��~y�������{|�=�Sh�=!?3}T��py�������db�9�lY��R�0��2��{����X T��`���Az�7�I)�]Ul'��΢�WgW�5.�E[��+����&?�jg�`��|�sL!k�O!�B�,�2zk��1�����C�'�%*KQ�2�[I�(l�)�j��~�f�)߸Ѵ(M��i*3kBn>_OH�F�Lv��ka9)��z~�n��j7r�`��[C�,��]�=,i�oK�����[M�U/AIM¸1Jz>�8��W�l�����-<]���ܗ"c+�Q�l�r[���`����3`�=˝ ����h8�1O��J<,��Ƽ"�֍$�$��n��4[s5�0�C��~�v6�Ɯ+��.�؟;/�zY�M[7���|/:[&-�E�=�Ψ��0&�E}�Z��(_O?�W����#�%E�'a��>������AdƑ�z���(Ml��}6�C R ��o�Q��rJ�=R�����]�	����!���=z��o�A�=�x$Jٴ����#� [�=��W��O�]i�u�4>����\Ц���K�!ދ��u�駮�9ď ��G>3�k�O��r�jT�Zy�f�w���U�)NЩ��MlX� 8�aԟ���{�O��k��v����+��*74�����6{{z}�mk�>)6b��M=�u�~�6���_�)]eǚ�C&;<n�k����6Y�r�$
��a�ㄙ�[jD�ڡ>Pu��h�����^s��Y��e�nX*/��V�+eWTm�և1N�?E25:Ģ�o�\9m�Q�S��C'sRwaq�P�y���&�kT{sU���3g���p�.�.:0:���"�l���.����~��i��T��:�#,(���*�l��F��~{�]t�+)l��O�� ����
��@/p1�;� y��/86%U0�!����	�9t��]>�?ڌ��+�*���?�I����3z�O�a��	�F�TS�P��qB��3WA�O�|X"��T�N"�}�r���[V�p�QG�5Ȟk�wG&� 6���T	��W��	�qw���s��?КF�a�����C\�`=|!�u�]f�(���|��Û�J>�iy�AV�i��/!G�+��֨����a��%��@Qj�|�U"/���	���w)y����?��l9,�_�PW�T��Q�\gV�4n���?q�Gy�2��(x����5��8��_^w%���S��l`eԳ�g�k�<;Z��R�W>�;�*tL�Tr&]�B�8�  ��vN�݁10�b� !<���	�k�1���&~IW���r6�PL�$!��o�m��؆n˳�"���__V�@*g��"e�MBNIؗ%l��FQ��hKZ�[
\@2��P�����Y�BΊ�F��y/��=ސ}{A��.���w� H^����J]�].�n�'����9O�	jr�@�U1o�g��+T�8p�)�w�M��[v�=�L���S匟����Ծn�[h�(Ps�IET��<Sd^�m��.��j�j6LU�{�6ZP��`��x<L2��X�Ֆݠ
q�F�)nv���Q_���>@I�̨{���3��֢� ���o���9D8�O?������$c�ZN|?���.i5]d����߬���+{����sBג3#M�9w�__��RF_ǌ��k�eR�:q͍��������$x$�|�#d��D��yw�X^���@6����8R�V�9��L`��K�n��sd�q��(�^��n��:%���s_k��
����X�?���D*�3��a����a,(�J�P =���h�Bm/��U�\�@-:���6�U�눂AY]���zUi*��p`TL㨁T�I����c���6�V~e)�	�Z�5g���<09l�R|�7=�f9�2���Vj��a�|?qZ���TUݞ�	�ط"Z �Y��JL��a3$�X��d�]����6i;���@[G�	��@$X��D�8,�Pb�tg%m�� p���}���`��+�գ:>��ݏ~�[����pa��י�C�b�ĳA������Tz n{L�����W�, VX��n�.�F�[��ra#�/Й7[�m��U�d�)|��	k���~_�Z�!�w#��������ѐ�!쥄��,bU�v�E0�1�}� /!����D��v��:N�j�aiQɻ�8�E�ӂ�q�2\�o�z�)s�~�)'G�v��P��n��">4��mB��XD�,��"͉���e���.�Qse����.g>)���1�
�>�~�q<2��Z	%<�""�&��u�4@�p���i�$JB��7�@�۷	�>b|��>O�]��R�����sd^����\��Ia͠�9Z7G��"�g*`�T[�@ �| h��OBq�u��A��.Y��<B�����[���v�̫�ك�9(o8({�1�h��y���~7�mƇg��S�[H�{�zN]8dM�����Y��P��Z-ZR�K��Rz�+��l�[6A���ݽ!�s�8�S���02�g���!%��g-��Һ1"j��M��*�P`L�6(l7������~u���ukN8�"�� Xd��e�i���tT�Y�&^�7�������<��cG��2��������M{Bn�5��/���	E�ƥTq\���hLh����%I�L�P�s�[� M=˳	8F+x.	��R �{�r������i)[z���@r7��$
_�$Z��>@�Q'��Oa�(��V�a��Ӻq���������U��םI���o�.r��Q�(� ��n���̳�T[*I�s����;J����`ۖ�R�e����W}m�����ڗQ�B������y���ˢ���L� ��.ύy�\Q��[�	qk�~ p��*f��\6�����^�n}v��f.��]�5P��;NDDf�:��e<��5�&ӆjR}�w�0&dԈW%lt�h;B��:!Q�5),���,���(�I7b������mw^���4�ǣ-y��<��Mn��Z�Ψ���f2��LD�m�Nڔ
^Q;�y��CO������6͖*�o�ޱ�Ry�'�8Prd��,�u.�:�9D�˾x1�+�ƸQ�Y����b��{�-|�BY.�Mfe����΂��$�R��ȱL�J;ז	2�p1�X�A%-�1?D� 3d&����Z�Ø��di�Cn�����Αb�-%��]=&c���%�u*�A���4/wz��M�A�4�l9@|�n	1�y>��%�w��cڧ�o���n���mX�-�@ﴕ���	��CEIm N+8�d���SU�H;�7��C|T�_+�`h?E���U�5����������*~��,$`_��2m�������	a1��nKF\�"�� ��Y�`5�����m�|��CȪH��#b�@O��?*����5D��5�$!ʹ���?�j}*�gl��]E�H�����K�Q+^o�hF�2՜G�d�g����}�v3cܓ�=��ƴi�D���\�݉U��ٷ�R��Wщ=�{5�$k�z�h���X���bC3�����{����ҋ�������VfhL��7�t���jE2z�='�z�:nY�	(�	��� ����tCZR晖=O���w�r��1��z{i��B���!1$?MY�	8V�>�=X�>
�)�`PEX����dR��|�#j/5wfܜ�M��N���N	ML����0�n5���+G��Ȍ�E&��n���/�]xM܅���!��3�U/��m��o>��	�tCۊU@��{��/T���Ue��T�\{�:�@LϨ j@��=qB>�/׬���<� ���iXBU��S�
���l�Yy7��I`M�UQ�h���pP$�5���b�ɮ���J"�ő=�s=�%H����!���K:J��f�Ȃ���x)�0i/?�t�@m�}i[8p:e����H�0c[�w#�2	w���R�O��?��5�A�~�~Ytm!#z�^̅�_���u�tQW�|�Vީ'u7!��R�=W����r+Nn#^�\��}��w
�X����
Uo@P��}�{����|�ӑ�Pc�V��v���X�����ⅷ��d���5�ӰP�'�����+t�ݲ�^՜ʰh�+��8�J��R�<��-���g��9�c�������R'h�����ܗ�pΒ��&]|nJjԝo�x5�I���[a�<�?}l"�M���N��F��	����mjZaUo���[�=E��l�Sk�0�dy�F����W;x���T���C�T�@�ߧ�5�������z��8�p�N��w��1�b-�3� Wr� F�Bk�nkWϱ0�u�d� r�g��R��<�@U(BRyE��͹k�$t驼
�-��[,-��eG�B�ϊ�p���"#�{]l��^�Tʙ�U�S�b��T�t`6[��7T$TMu���4��=
�j�x��(���b$d��\2�_�C8f�J�R�7^K2t������x�o^����rp�֏��A��1[6��_�
f�l?1�6.M~|Hm�&���Տ9��n�_����LZ^?Yo�(��i���Y��+�!����\zY*�����0IJ��J8��9`ϮG��cG�����{Z�E�ZW/���B��K��a��-1}C��D��ےqv�S� ��A<�d�7�ێ���� E���F��͉\������!�K���X�*�����t���9��L�����<|���v#i�[f�a��儰��c�=���������4Dg�:���h�>eˢbk�jQl𬤻2��.[���(�ݨDtt�%n��O�N��j΃Ձu3JÚ��b*�./��zr_������=�d�!O��� ��k��Źʯs��Y�T`<Q���xGL��
�r��8��S�[�-���>�W�Ÿx���衪*��� {n�^�wsO_ʮ������,:X���?��i�`8)L]7j��%�Bt8�c�mwo-ۍe�<Uy��e�;۫�:M��?Wp	��R�	�~~����7���d6O��Ȓ�Ը󣇈y@5�i�X��t�=CȀ�=<���}{j���*!q
�~���pf�L�.?ޘqB �VmrP"�҄���aY�?��̿sp��H��K�Ll����((ix��\�V��]�nV���1��葚0by'l�!L���S4���
� ,�p���HA�*�^ZS_�ND�X��{�C����7kUhs��ڨ���'T8an��q�!�����.ގ��Ow��lj{�eѩS�X����Tt��rĐ7['�5u<Mz���\��y��J��z�����
�I��z)v�K٫��ɓ� ���RL?W�� �I�]�yBh��v�gG'�:g��iw�K�Z��N�Ƽ�R�pof_����1��!6@~`�%T��~�}h�":CRA(�u�.2��D1�!��`m$2X�:�
��]����6��5�X�k䒗����Cy��r��P�Z��Fcl�zH3�#�<Ş�ʈ��T�Y�ꏧ鵞>p�y���^�mO�e��,A#����&#K�uMD~{�7�rr� ?�Cas��?�~���	�7,	rށa(ȫЉ6�в�U�� g��]���}C`$~!4uQ����J��Hë��Ii@w�rW/��T����U>��}X�=�-'dN��-kPT�n�Fײ%S���(l�p�]|=f�H҅�����m�.Xy���cqveA�]���i+���H�x큡Y��(�eT�z��̈́_�1H��+07=U�
��"��/�&'ፓI���,~y��ᣢ���|kh��EJ	���=5hL���rfh���"�Y�h���fPh�v��&ӧ&���ܞ��U ��/�>ݍ\:�˪��9�v�$tU�4,�C�`_�7,`~���F�x݈��H#���p��x?���v��|ʟ�W�F�������N�:S�zo�#�l�=KBl��F�N������AG���^:��_�K�˛
�=K�::�����H$��P��Q�����c&��ŎO�9�,�&/Ȳ�"����i������N�Яc��7}����t�R~[8[o�"mE۰ӯ�F]���M��"�S㔶�5�$���k��T^peF��l�a0 �f�	r4��8Dj8ʴ�⚫�߫͵�` ��K�t���N��I��(�\���F�*s�g�5u҃�,$TR���X/G$M^��O����*�F-�o�I�o.����P�2L�[Q�G����O5�b�%����hl�y5����Rf�
7�t��jT�0h��b�`��7�����맵s�t�҄B��;k7�m�}ğ��m��p��tR��݇��t�2~� �I J�A���C��j��xq���Z�O^�a?�7�h�O�l��HjO��&Lx��Pr=�-����V
�.�0����珵�d:��Lv!�S��^N�#���CT���J:�(�/dI�6M�;Ts�蘤ܷ�ў��mf{�W����1���˯�i�i�F��9��Kl�ӸhϧG$ֲtSf�3�(��Ƅ_�u�޹�ܛ�_�'2J)~�/gU{ɰ��M*�������~�����ӗl�e�����d�O^�-f>���|�ൔzr?o1��|=0�~���6�쏻�����Oi��	Zn�8Q�wp�^�N~䧻4~u1mA	�C�mcT@V��tHf��s0�5����^���ܾ��ti����B��Y��u=��q2��<�C�>h |)
���\ɿMF}ZD��S�;��U��h�!���>��P�$��U��*�lضو���b��a3w��0џ�<: 6�(�v�$7V��-"�ɑqа�S����a[2���Ϩ��G8�ax��1� �ֻcE������/�
�wV�NEyO^[3��@OZ��+F�	�5�Cx{�p����2z&1g-��#퀛���!�+��m#���cͦ�;�mk6��Ū�`�f�h �mܸs+�J��t!�I����2��Y�/Գꇲ�<��@�h�5:G�h�50H��[�\�5�_�ߘP�T�I��t�1��\/6e��9)#]�!:E��a.�I���}ẑ����YB#�M�&J�����t�ÖY�F_�WM�����f���x�A�V�Nw
�6j�|��d�?����eY����Q��'@�h+��I��<�� ��/�ZS��U"��� *��7�9��wт��ͨ���x��G�yPv�Z�)�Td��Q�t��M�"3[L!R�R��m\����݌�-[}��(v�W�WKd��7t��5	P�:���,�����4D�p6�,�W�Z����	'g��X����d9�,�if�ۧ\�����H빞ES� );�k�o/�Tjz��>�?���1(Dh%�� ?�D�b��ο8�B���kG�^K�e[�Ó��uM��:��z�EqQ�J&�mH}�9�`O�'�ڑ��g?�(�yAΈL���J�Ԃ��a/)�3�+��<ĳ��	n9���&7k�#d�ê-֓ 
��jV�2�zO�����/�O�hæ�.��5�p]�ѷ�1)RN�m܎2�5h��������M��'6�e���60��	�Ǔx��y�d^�/��0�^��	�V@��#qՋ�hk�5�g��Cn�
���z	j��S��WH�D��h���<.u`����B%g}6���i\�;��3�i��Ы�,g�s�[���z����$��4w0��C��m�'�g������=���fu/�eK��9���Ֆ]���D��\�z�l�W�19��,
��/ʘT�L�5�ڔ~�Q����Ln&��fЄ�+�/c�Z��Щ�aS�f[�Y�ywe"�(�����_����4X~ ����&��t\����=��h���Y蒴�H����#7�A�K�R�:��)%���ۍ8|���F��'5$�#��#}f��=�M�����8{(��5k.����� �3�b�n�}gz������0�
P}D?��8�����	*_2�c�Ƒ�\��o��S! ���Cem����!�87|`Pk�$��y1����4�"��Y�����.�W���ӱ�s�a�.ց��� ��(:y;!5�9�Ll��$W#4�	u��8&u�9�`;A+*���?� �����.����&w����$	���6�;:Ƞi?RI����7t�/�A����J�Z��M��=��N���YN99�Z�z�&e�Y�y;v#8�!O4�)��OLf��v삀�Qڠ�-'�"��.7"��s�]����V����3����5*57�i֌߅z�mdzʄ�W���ɒ��
<�ָo�c{K���{�ݘ&cVy���Q��B2���'&�ֺ��LX�	̷�?c��&QJ�67�mM�*�`y�8��0β�tfY��ZW�u�[ꚟp#��%Q�\׹�p{-#�`��:�u������'�F�F��,��B��3Н�vT[z�}Z�$�1��՝p�bd�)�rTb%��O��@�0���/�#I���B��̈G^�R�Ւ3ܭ(��E{T ״�4{	���H�^��p[ 4
�-��l�}uC8�L�Q�i�����õ��a�⚩>r���q��N=eh�&���Ź�u���Ys��`���lz���4%�m���@��%H)lc��#�e'��3�ĳ�H�V��0�M����������=�{l�o��,3��H�����b��^ޟ���N����F7D���.S���$0�;�3`O�ʏ��XT�����s���(��k��g%:�WXU�!��>n��5��]��]P��:r_2��c���?T��]a���hcЧ���NE�E�fLt�Г���j�M��Հ5�	�V)��1u5F��rv@rQg7�Y�5��bl��$$��Y�I99���H�'R������n���-��tЈ?��R��*�F�l6uNN��{0`S��'�+���#���kV����g���)��	�%��g9��Fm(�@��Nc}�U���5&A���|�ƪc�@ī�;��d?]F������m�� �+
>HX��a�,�8�������f�C�"��즥���/'0!�XlR0�9�d��ʗڰ��%�[a�+�г���0�񑿰-B9���w�g�Ҫ	�
��P�K�g�KoL�]uK�'���'�W�]��.��,4��Ω7�N2Nj)R
iD;tq�ҟ�%�aW3r	Z0��BG�S�Y>��Zៀt#�r��<�v���+ܮ5� �6�ST��c'���Ix�5�7�5�Y��1�J�z�d�)|��*�$Vh\��]�  v�C:����Q�LL�������Yc��m;�6��"Y]�k�-%|�]"0�,�$?�+�4�٠��%r��c�a/3�n�R~8�����ƃ�d�VG����:��!���i�P��*���XG��r���n��Q�Z>������_���aA)s�8}����h�I��O��YX��������," �8K��ڷ���kй�Ex�w�o\���^,�
=�|]���H������.��I�����y%4wCD���Ή��\�҉=6˞��r���!��}/i��BJY'����DG��Sӹ������D#��� C5�+�$S�l����ƋYB,.6몷�~�)������5��P0���{:Nhr)���P�a�u4M�̊?Q�6S��:��A&oَ�K6'I��R�`P�c֤.��/}z��_(��{���F3������E���BW �l{@�E��*��)ĉwmH߭�ف!-�;�D5ժ���9�����`�hf=o�I�����t
bH�M�_#/�r�U��ߕ�v���Mr���(b�|�Pq�*fsn�}�k�8L�.˵�z���N���e�MM�. h���ZI�b�?"�Z��:m�8��Ȩ[��վ�j�yz��&e�֕RF�	6��'��z�JT��كx+&4߰���{d�3�?n��
jyr�0|����	vn�Η�n?�	���#|(q��09P���l<[�.��~-�,*.���p�R�*�0o�N�u�:�k��>�� HD��~V[`"�ء����y����O�?�_�"��h�fS�����Ϧ��!������{����]S��Τ���~�)���=�Q	9gK�#��=�y���ގ���Aո��H��lo����ޥ��DO�o�A���N����iQ8��:P8/������@
Isr����;�s��okO�}��V$XE�i�=c��ޗ�-w ?�5Q�#ZԄԸ	����V�^N�^p��<iʀyd
�`�J5�,�DklSvִi��f���;� ����>X�G�j@��g��yd���s��S��ʸ����e.�뱀-�Z`���"uG\�WCt3v���-a��:q��=�WY	.'*6Y�m칵��ԸC�#�]I]s�et�buJ���Ƥ��7�b,m|�j�أ�Y�<`��leC�:}���k�L�����|�Μ18ӈ��$���q�J�fez^ˊ��:��]�1_bJ-B�ڵI�+bC�,R[�Uɠ�#�d3k8�G�D����i�"�F�]��L��M+BJj]x(V�d�>��󨟻��/�vJ���	���[(�n�����QH�p�[�I&i�U|a����ٲg;��h���ז�C�F[�wt2�/�՝!D���N��w�z�+�3Z�m
��UN[��k9J��+#(�j-we+l�J��$���1�7��DA=�5��H[P���a�Ϧ�.GK�� }�]��x��J��#(����Ս�'7N�P�}����l, r9�b����4A[��a�5�r�6�����l�df�(��&&!6�^�.�j��S���HL�r��S�Y��<7�Mؠ�^
��������(�F�$:�u<HRȐ�ݛ��6�=)[�m�p��7��5�C���RA�#��wf�w��}L��q���K�T�.�N�=�}�_�I��Ɏ#3���ڌD��>h.Bq��竡'��c+��!���"2Ģ�0o��/9�*��WR��d"W�x�}��=��Ȱ��a�/��@���GE�jA�/LE5��(G����q�ơ[�&ʧ�k�$t��,��z��"�:1�����?z�����L#n�O���k����6�W4}��M��K�E�˵wD^�~������Q�d6�g�mz�{b��J��zQ������0��V��ۗ�)e�ӽ@���]D2y��8ﮂ;?4h�N��NB<��)�ŒQ�@�~P�іx҆�5��7{��l"�8�3���%CPh��iB��3W2hu���3>Z2�ľcH�_�vЯ��Ց��^��(�ח-�L:*��>rӣ��G#����o��z�h�ݧ���(���~>�=��w��V�*q����?f����\��ɰe�
%`����V�m�F�	�S�Mj�󍠖l6*�۪F�Ưw�c��<�kYVg�g;��[* �At'��r�����Xj���H��]���i��-^4�,� ��'�V�R�Vg)P�&�?l�@L�j2Z��v�b�����4ڤ��:��1�=8�?�Ep��2�r����O^��8��q_���;b�9�c��]fQ_q�:����ۺn�-��C������ ���3���˭�uF��/�M5�J�kgK[&���S��c-��VV�H�+��i�ybQԜ�$-�<�S1Ӛ+8��B��a� So�y�#W�)�ºiҤ�,a���oW��� R������̈c=L�dS�a�����͟�2�P;�<
��S:.̨q���V��CPZ='*���´ز�Ex$��ߋ���4�c�f��z���I��C��y����$�y��*P^�E{��Z��/U�x rTh?Qi����Z���8��n���b����@Z����j�	�K�T?�&��\��?�z"qo���UT!|2����!9ر}\V�&��>��~Y)�/$����f�����	ĸ�^�"�_@�rG���?�'ϰ��v���2�Vp�{���Y4���skn����\>
")VҶ�	j��j/$�m�~R�����w]�Ǖߗ��רN�0��qF��N�~]$/Z|};��*���^C��.�{�0�ߙR/7z^���20^��X����M��"�����wl
�}E0^Y*Ta�ݡ�v�=�� ��,C�}kяP�f}gH.i[.E�\���oR�J��@+���@3��<r]�¹�Ϊh�"R	iKa�[�D�!�"J���J-׬�ǨC�C�EٶJn�76�<��x���/5m��crRy�=�[ee�
���Efp��-iv(�U2�7� �Ά[c�@�����z!�Ip��K�OS�z�]w�8����}k�d��l
)�����U̮�"G��E���; �g����J�T���#x���G(�z\���&kCj���`�3|+J�ύS����g<�aU�X����d2)����*q�6�h������i~����#�����7��C�����a)צ�k}�5<>g�%����=-�t)���8�5�)s;q�ڒ
;���r�D*A.��|mY�|�1а}�O�/����Q9]�u%"���j4�9#3��p^Ύ0\�&��Ug��H~�*�9h�PǍ�yw�+[�2��b6�%D2��+V�b�םsd�jL���XPO�BA���
��V,��v2.8��������Dr�<&�wʝ�j��W��H�a`�8g"���[ĵc�1���M��S�x�
h���A����B{�>`��T@LS��V�ΜꟘ|:�N��^�y%xm�88���V����>m�S���������g�*!ʿ���"|����z�{�Iq����$k���UуQ}s�� 'V&=M��T�<�B1�OP���{f6<��9���rѽb��`a֞�~��{p_��e�1�3�D5��KT	���S��y�;�Í��*�ճBP���b�wTXpL��Lo�ݩ�p��-v�m���g���2���֥�$AZ�Q6���z�)0�5)�2p�;��]��P��&S�}m֤�F�(��.b[���R�|��Ջ�4���n��:� ˁ�3y/0w��7x��P" v�/�S����܌n��ΪֻM� ͽ>W�L���b`��:���0G]M�#B�tl*�1�װ;�$�l����uK6)���9��[0��1PQ:����$Y����׿�47w-���x|(�۩����t�bjb����:�fKGi�����L��7I���,�EpQ��O��IK�a"�b�g�	�b|jL�u
H���,j�$��#U�5��B?{@�,�R�=�&)�R�+L�B��h�9�U	���9u�>�;��(�����������k��?��.�~~�a��p#��z�A@-'�S�3ȟ����V��N��Wy�>F�ʓ�ظ��י}����+70+�@���y$�9+ �Dp�-���[��;Q�Iy.:;o�8�J��9]U���]�cdZ7��B\~g*������T��b�Qjt<⎱$�]��n��%T���$����ѿ��}�H���:���:� �/ΎC�8J6d2��>����L���������YT��-��	�~$,S�7��z�j7�N�RA���J����Ghp����� �!ےxYvrY��Bϻ
���0�@Ɋ��H۞�<|�����uu�u�%I�b�X����x,m�V��e�2��K[�4�CG������
����pu4�4�Z��e:[��ŰQ봈'X
AjWX�o��@f�
WO^�Q�E�sr�\�9(4�W+A~��ËڎM�`?�7��,�S�^QR��qB9E��>5��}�A�p,I�m���1o��dcj����������#���$�aP}��%Q�5N�&�zY.�Dم�Ae?��:�6}�H����:b1�[�~ϭ`0�5���'�@�#�Dt�7�c�˱���38�y�#n�|Sf@Li%R�Į�I�&
�\�a@����ٴ3
�\b#׌���R?mmr�V�x�9Q�m
AjV\7��b����'�h������t���<���"|P���ʻ?\�Sl>M���β�`� dzwT��qL#�������x[���v^��S�Fs�-7I�^�	MN�d���������}�~��<�#���k��J.��\ʬ�2�e�G������λM�J� G6��PY��1 �h��|T��IO�>�j���o�����(�<�����?䅖�J잴��c�B���(�*��R6�=8���.�ͳ&>:��ݩ��S��x���4��w"����#�:U��	��% ����6NM&	��S˗+C)�y�s.�]/��2��=�`!�5X���B�8[�ڰ�����Ft���~Ea*���*_��h�0g�T��1~���U[e��8>�kn��=�-�$�Wp��3�?)�^��&e�I��M���w獵5T{�E�������t�a�ܬRq���V�F�� #
L��@O��	�IBu�_ї�\'��Qyk��"T;\�<�EQN#k��p7ⲵ� �5�B2����%V��{H��m�!�e!�C߰�58�MW��kXI[.�;��9�+��@��L���[Pܦ��"��saܯZ�bf谹1�+��q�A6��U�hlοp�	y`Z
�:����#w�ÚFσ9=��!Lءx�H/�F���>\�Pz����yb� �:qF�z���vڐ��OJle Nn�N���*�����Py`pZ%@�h!	�����6MpG�Y�,@ �h�
)�Q�9�}y7Z�m|�㧉�Etܜ;�  ��E[�Y3����vu�`����@�B�H�ƠqD&���W���ᬸ�_1to�MlG���m�/�Ϊj����#���/z	|�,���2_U���5��lR)�Ь�őө���-
���AF��	I��"�f�:��v��,,��3�;޽*`5��sz[DX|cH`/ﴅsPR�=CwN>�}Nİ��	��j���1#E꿝J�A ݝ�zh|8P��"�L��f����H�	[�>�R/GD��ͫ&v���I��U����錭QŰ� �6�Gkt���z�I����1�{���4�,��iP�e�� O��;�7���L3�����e#��o�ʴ���u���K8b%cR��_�4�}�vw&�Ѣ'�Ft�_���8B|s���j�e��Tp���>��E�.��[��L��񼏄+c�S����;�z�Yd��G��kr�����GXr�5��}&)��rf��U�m�`5w������ş��ҡ�={�#��c1?6#�] ����Y���'k���6�w�ߕW0[���0�sC��z4=�Hx�}��Ӡ!�"ݷ��Ѥ�H�h�=��V�{'��Íc�g��d�E��ȵ��7��N�@�(�UL��I���1v�1�����K���%��@�ꖡ�{%��M@��v� ��t[�i����
�n#���KO�CIeD�`��x�j¥
���"c$P�K�9]%	�'���X�$�[��XZP��$�=��j-�7��h����n|>�յ�.��p:	��4^��8�>�[lP���(�B��]ZF����x臃���QnΙX�C~P�6/!��V�a�����;�tŜ߃�ni����a"���ǳr�Y	��E=mh٣K4P��dn�hm����ӗ�����ծ5.r2:�U��\�E���@qdHR����H����9�;�4H�$��0���F~��qx�7�O@�p�#�'�d��pU2�PR����e��b���3����4�8�+�#��������~�%?�z��(�����IK�E�Nې�g01���
� �J�����}�P�rR������I#-	�+4O�V-!�4��
[ٝ��4&�c��R�8w���jS����{q�ǮU��F��ۉ��I�÷M� ���0���T�����ÜZ���G��6�J�A�z	���{ л��쪩��;#�0��כ~���2t�X����pU�hϻ]�j�������Hb=�%���QU�ʰ���2'U�Qe�x���� �k�e?�w�i�*������ZO������ީ�����4��S]��E���3�/��F��S:����{�T�3��kT�/��/�i�"�����ު��)M��·D=�ٵѵ�W���!� ��������H[CG��K_�嫑[� �SI�Te�������1+J��N�0����C3�)��=&�kQ+'��x�V�Τe{�+;��|���ٷ 6D��2�n}�n띄���mf���&�ќ�r-El�wrh1e�N�.�ՙ+q�4g�T�8TI��/�Q�� �݆����� :�4���[,�`Ԉ��rQ���]��F6��Y9B�I�%�4(z��F�9�2O���B#�m��͉��>b]ґ2� d�c$���I���*~J�p��|�h�m�?�o+J�拧�+86U�<!r��5���j]Dg�h@@�Ws�0���0H�p��(�����fTe6d��7P��	*��9�1��V�3�����X�*0IU���%�\��0_:|:��+��Zu�}���4��˞NC��;��wo�H�`�?��ܨ����"��0��0� b�T�]�2?#�5�s�%(ٻR
��禳Q���Cw�_�Y����$N-����e����R=x=:�&�3�o#��VS��5���} G�Q�t�k�Ҧ}1:����69a �d���Ǐ��r�n��.����.I��e���� �-�qE~���Np�o�ݱӑm-�����!�h��E0�Ҫ��8a-q8���g�t9H߷���W��)@#]&_�ă�"�z��H���Zd��t�i��q�j�� 蜄G���x��x�j�ް}Uq�ucϔ�����u�õ	�z˹e_K�yc�C�nGT���\�WDįY%�u7�ː1�����������ɻG�kd��������k��[�çR�$5�=&�͉�Z D�T�uL#_F�z�w�m5�8ͅ�O�J7�[��m,��!��BVyN2�TlV���U��	p Ӿ�<����M�B�F�����5		�b�����[,8p�+�6��+�k�T>��!\J9RL	�QI,1l��j�Ʃc��+^���ٲM��H�Z��8��\��������19��<sM9o�c��gzl/��1x���Y�E*��������X#�ú�_�ڮ �:�:�uX�
Y���M�����	��Hs.�E��k]��j���A����G֑g�v�P׺�t��+r�8U
�}�ȇm�ߵ��
=`����T����h����DN���Sa���b(�&��	��l��U�[��8��K*V�;5�[�@����/��8@�y3#V��a�wɲ@�ʉƠ��L�\�x��Z2�&Ps�Ks�w|���ڟ*���¶�fja��XXb��6f�1Yz�vK0��������`�]O0����r?�-�l1�\&s�����9��dp���1��j_��U>ޛ�f�̖�}~f?��NN�J�&�5v&YY�km�����y<U2��jC�J��o���bI�,.,b{�\�*�}�'����\V1ћ��tz�F��M���#��x߹@�9�9pa�r��9>��v7�֯�3fo����1��@����Ɏ>�"-�5-"ϧP3{ŹS3�r F�;��q�t~^�+��R��	���@�t�<mg]�sNV�]�2�pKK��g����R6��'�|P�� $���g�w0z.�	V����o`�����].�����"�F�>����-=~ɥ^Eq!��$0/���B����,��?��0JZ��g��t��b��˳�Z'�5pu�'�
-�䶪 ��6Zy`�Q��\)@`�/���<O�U'T�����������֪N	�����H����ЩoAm�-�3B�����e�[8��ơA<sJ�g_� �U1Z�p⿋���rק ��^�̗�F��+����o�&AS<�����?=<��l��W��>�V(x˭�P3�7��{�o7���yg���D� t�T�"�c�F���\�>*�U�����W�J�bV8�~�X�7�8V��v6�M���d4AL=�;AG\qU�����)f�iX��Տ�x��1ak(��U⣐ 99I p�mLPs6��8�З(њ�(&�ի�ŏ�q�̭]`n���@�6/ưÃ{�O*�[�b�+��v#����p�lʫ�o0Z^�1F�0Ji��TҞ絞sۣ�8������NKxu4���a �\��[���������8�)1�k�g�ĥ�����6?F����e�5j��Ƌ��|�1
��剧ZPY�|�m�s�/[Wv��Y`�}�2�`A��5�Y��3�g�j<<JE�`f�>�8�s�?�������[��/ш������}����D�z��e~�؏Y��Ʊ݈�DĞ�����q��	�W)�w-�/C���
i!�m���k��y�������BJ-�:����*P�d�f�#m�q=��ޒ����Y?���&�����q�xc?���^�v����9���	}����X/]{B��f�L@�Ēu����Mژa����F�̐�6&��ν�|/.+�$Y�폁8t��B��:���+���ɓAĲ�j{RU��B��:�ȩ�GG����!/I^&�#i	�u�Xd f���z�E��^8��y�-
-����Lԧ�����Nd������9	� vN�]i�hn�q
�0xEdW�?��)b!\ʿ��b��}Q�1r�E.t�&M��b@.���꬞^�O�}���+�+xQ�!E����\�xrZ�i��7����� ��/@�键}�e}� ߌ5��C<ރ��g��L3�bL�U��\�R���en˹?����N��}�k��	�S�=9[a��Ek�|�ф߸D�\dg� �fXO U��Z
&�4\0�Ǎ�[�۸����g0����82��w�F��lPz3�%�C���{z�Z��	P(!o>(��1�e��l�DZns򆮷ǹq�������W�V��{]�~SX������h�{�/�e�<�]l1�1�|�K5%�m݊�,�I�q�j��Ǧp�s�8��{�ը&'�*l�Ɨ/E��<�+Uf��>L��Z!���F�֎+|Nd�i<{�֥qO!F-��W�Z�"ј�K�j>�6ۼ�Qܩ�xq��UI��Ke���P�Ǌ�h&��d�f�S.ⳑ��Q��pNp�9(���`�I앝�hN���t�p��RL@��� OU�K�c�w���Ƹ����Ϲ2�Œ�A��ƅ��~��Y�����?m��%!��H��		/�ۡ] 6N_,��k�~���4�7���aI�:
�:�	��,�n�#9d��/��̆ )G�A0�G�F(wJ �B��Xf��4��m��m��ي�9�p&�z2Xy����T��Cg���"��h�8���c��5�-mM��;�I�
1�s ���BH�x�������O"��yӜx
��xZ�7 P��%�����":�PU�n +�$���h�&n������u.�wp�?2�ȡPV�0�b|�rG�ź$\�H��(k�w�񪳜��4)~"��z��TIh^/����#�t�:���t~���,M>�ض.|��_	�N=�4.x���%�3yv��
����}�W�B����~�(pt���=w�ݹ����σqm����H����Kܰ��/�D�6{�w����胔�2���?H1S:�Z�2z�˨FW��mG��@�K��0orT0�c�@�r���p9ݑI_��0��:�AqU�\�$�2g��]�p)2��m�LI#��WZ��`Q&m�)0�7y��?����7~�{x�R5�L�|^��4� Ƶ8��;�~JBƶ�*�{2�p��y��F�����,�����!�����f-KY�6����+1�a�D
�{vԝYX�!�t����n�Q�!���͖�ZS�����.W1���[���N����73 �\ڠ����#��z0���JUA}bɸk����ޅOMJ��, ��:�������3B%V����F6	mH�!{ȗ2���+�� �A�[��dqa�M�%��it�C�"��?���	���C���S�i�WqnI_��ݏՊ�o�~0�;��� 㔨�=m!hQj%�PjN���=[��������i{�ۀ�sY�����`�iaϺ����e��b�/J�KW���qAȼ#����q���T�'_tNZȖ�j�{�0��힡�n�3c�D�C!�D�vo^X���/�n��7`���w�â�������Vu#8��r[�f��A�l�)Y�������/c�!��ЋU7A�`�Ҧ��wo-�6LF6 8�%� �	�1�q
0�H`�*�R�����驩;�QcV���#?muI�bF�+[E���d��������rӷ�i)N�:�6_�����";���
SSdI7^�`�<����5����'����@��L`��A���� 8��5u��"�O"��uL���=&���)�i=aT�\��#}Jsz��6%��p,gL:Ly B�e*��j�ƙ�#��=-�-��I'@p1X82T�}J>�M�_A���6��jX�o�JO�׽`�Ds���$P�.��v�W-�t?]�#W�a�d�z<ݪ������SGt$m���^@%Δ
�q<��J�W�$��[<&��V [�r��E�d���w�l� L�6�v�)�i�XO�Sl��q�����ʊ)��i�$�&��B��o�^馞7�M�^8�m$!�����`VM�#̿/b-�A��fkJ���	(�����><��>�w�y�cvb����6L�$K�'Pg��={����l�`�"U��rmr;�&}�r����oh�xޑ'K���=�o�GWX���K��6�x�ar7��(���兘`,mL��4q߹;�M�Ӂ��uJg�4�fZ�� �s�8h�n��=Y}-w"������:�4��]_�H�M&���c�S�%O�D�[Q����ƻ�� ʬt:���T#�qh�o���w���5���v(O�rt��-G?M���$w�`��6W�ú��^ӝ|���
k�Ҩ��P�Ef���r2ߓ���y�yj�w�.���tЭ�F;��|_�d��N��Vf)���?.;N+RM!&����O
�6��AA�o��n6)���ڸc�[+�(�	��j���#k�v)�ن�Zϣ���9ZZm;�˞OƞO#��SS]��Ll0�~T��!*L�)qJ]U�Q���s[��.8�yJR�dL �>���_����T9J�/�������pL��x�)_�Oy�
��n�A��!|����!˰Z��ְ{�&"�n�@a������6w�vO]��LdrX��P I�t«�=���/�it;�J�����3HH�T,�AfP~�=������6�%^��b�w"�
�ZM �˺E��N���@	����9d��C�f�<�6�M)&�V9d���V�����h��㇍D}�	P����(��Mo;����bL���/�����/�2�t�`f)�������5`�}���b��7@�@x�:NR�ݿ~��BC�{�ڂ�~0lr Rg.ɑOo��E��K_[�a.��7��2Z�:nҕ4�3|��>Y�bH��<�\6FI�]�F���%��\w�qP�lL����o�`L5����P+�A ���5h�b:s	M^򦭂�5G9:]�4��������PU'y��?���7�M�@8vz���7g~ˈ�'�T���v#���҂��$�.ϒ��^���7]��a�&c��%MGW�.�d�6J�8`��Н�LMۦ��˗X�!ޟ���O��S�V�F�DB:�ٔ��c��˼��%���x���jO#쥗�����X|:�f����]Y�X���D��MY�PB��\?�m�N!-b�$�:�)xf�B��/��Z���pa_�e u��Ù	J��]�:{��3�┽n�ٹ!�&����.)��>.X^���6nW%d���b���갎�rQ>
sC�W�?�#Va�:�r�#��p���spf�r����w���.�&]���uT���Ûvlm~JC�@(�"�  ��B��5J\'s	6L��s;D���Y�֑@8��)٦a��L��'e S��'L֎�Z=�舆 ��>j4���?��z(al�_-�j��t�V�[9��*|��Y���}���;i�ǒG"�)��'���>У���y�o3>}��\4uH��^�<����?"!)�69��E%_��pf��jH�-kY|F`JL6��9v�9坔}P��_�v���?O�l �sM.-�vJaա��X��I�6�$�x-M�>����	�7=FB���Z�0C\w�����q��U;4v�Zk����H;I��|�T0����<"^h��*j��wˁE'�U��?hծUHx����8�<���~�IYh���Ј�[}�5�`(�!�Cb>���/ٳ�7b:�3�T#2+T����iRm��#޼:'���U׼���$T����TA���@�tA#dT!!���`������A��$�3g��.'.���I�����-�>�%Ȥ���Ny�v��b�)h �pm�y(H�ވ|��}J�s|�/��e��+uI8�O|;�S�5k�$�	\f�w�{J��8�KM;䪦����ݦpQB+�� a�Q-����Y��P 3鹰���;ۼRF(\�r�<;��ϓ��g#P�<n�6��VDRI��ரc��tvbES7~��.��Ý�%�l8*0���`�+�ӫH�
V/LL�c�H�u�GY����oT�lʄnΘ
��F�-�X�߿��ނ�f������ۿ��,t�&�Z�S�.Z]��3��ܗ�`�Q�2�����<+� ��!4�ۏK���6��~~d��J�cwQ����iz6�����!Yď�sJc��_�s'*��q���/�T�9�hd����)kdP7¾�}n�1�}j#�a�-�r���5�z�w�rߥy�D^pi�ְԿx*G��d~��T� �B�`��������Cbǔ�'�O����M��]���2 lԫ\ހ�� ]ƻ.	u�)b�ъF�|�M�J��E'g�A�*Ȥ��B@��׮��jϣV��.�ܬ�����P�q&}D�L�д8���,�3�-��DP�B�y��Q����1�7e��ԋ����cE�7ܫw�I�1���q�����E��43E��r��W��F��2ό,���]���=d0��Y��>���r���/e��\Cm��z�^������qP2�$��h�+�\�Y4��vѐ�|�{�*�쇅O�N��>�#����@��\!,�=ˬ92.�Ǉ���Ǳ2!��!�Fs�X(<�1��KXk�����C%����l�K��/2b}�=V�Br�-�k0�t2؇��]o4��h�؊ݍ��7 
��,�k�����~�WZ�u"v�3���m�%v`EC9s`?�4G�|ʭ2n�r ssOØ��j�$h�h}�QEw�A����÷�:ҳƀ��=�m%XX��\P���Z�}g�Gw���v��=!4-���↑r�}�>h��6u sH{&+^$|����L%P�~��俩`�~��@=��m�
'���,���O
��]y��L�&��e��Vz�XN�d9J(�X�$LA��g�v�4�J��H�1�����\s.b����'Q�a����o� .i�Ϭ�UR\dY���f��Ղ�q?�I��
Y(���0)I��N�::�{ѱ�)���	<��\���2̸K-i��q�f��?�
��iF�7���J?���=_W��	��$l�|���������K�5�S���:,u%"�Twr������?%�� A$\E�{�Xo|��ز>�~�#e�s�x�2Y��p��ϓua| �m��%`.�H�b����K�~l�+
�,�6��]������C<��X ��ɕm}��%+@�[ЅǔNt�}ݱJ��׏��a���v��v�y�	���^��ʚ���0哯X#	�gbeEIL�PrQʺ0�g��=a��)�I�3�M�E���|H�Z���|9����+��о	RC"4>f�G������s�q�b OAX�s	|z�����A-*�4�Z�=TQ:��e��0�}���=V�T�9��Uv�RƭPY]��i��%G{��X^���?<�-M�����P�?��A<���6�E�M�J�Jէ�
D�f����j|�=k�	2L��닡��`NP�&��M���ox��Ӫ8�t��J��u^�fȌ|��P%<	��^���m@��j=EюjTR�J�S�7,��c���dUg��|<�l� Xx���'>G��H /|�`Ȅ�{ï�����Nhի��BL�h4w�7w�����Z�`-�Z��z��z+pCr+��2��D�Q���e�GnV�Ⳕ+���0�y�-w��R�[���0�ξl�z�!3���Č�ՎA�v~���2CЪt����5�rT��l���W��*�W
�AxQ矧 `C�fe`���\�q�ƙ��|��s�νP���}�/��Q��m�&s��V��`!̰�ٌ��y�=u'�K$��D?u���0�in����B������]��MSqH�e�����vM��C�=E��D^F� 3��/�l��!Q	29eBkqOv�i�yh�2G�t�XR��Q	z��a5��T�CAE��keڅ��Z�13z�!!wŰ�8�4 �U �H\��{�X��qO���)&�X!�"���v7iIV�ë:)�Н�F�<�����)�n�"�q�����ɓ�a�wٻ���3�|h�ҧt$<&����Eڻ�wfX�[�^����__de�`���C�Ͷ�m�(Joh`3�3�{q�I�Ay��	M��8%�(B��:��L����k����1C���T�P�"W�@�K����2[<�����6V�׀kv/P3��+�@*c����������2#j���xT�W[mjV��K(���Q��PtR�-+S$�F����9BC�(^��bDȌ[cKV<S��]ɂ��Q�k�����~���/íg���#�����ӕsn�^=�?�?��1z�I�ʭ&�u�1�K�F���E�!I�� K�j���?wOsp1�_��g��ڪw�5��7�\ݰ"����o�&|�Dpd�(5RG�!O����\�<����w�&�� x�7/���à��Z-�������_�m���i�w%^����7�⒊c�xUH� Uh|-1��)�!G��gfWrm��;g}���J-,��\/w�YQ��O��GQ�1�:��+ ��P.Ch�;�S���Y��PrY7�!�[
f��ޡ\�X������v����g�,r�6�������3ZB1����論�<�=�P�,����Sp2\���z>�g�~��e���/Zz���q*1�z�����U`�̾�Y���J�橎�6k����Y	(
bjq���~X�z@���MM
��%�ڿh�bC�ǜ��K��-qR���H浙�8�\����}=�{,Ox��?We�~��՟�ȽݥN��כLܩ�pM�9m�b˹/��?^�]��a���/�+�\tE����M\><���#����Y��td �<B���-k���I$E��n��s��_�g�7������uH�lbQS�Q|RƱ�l�X)Q��O�����.3�\���,]�cU����N�4���wy�HӾ���3�J�W�^w� ���N�G���mX��nL��a]sK�o�(|*�|+�-��VTJ/g�)�Z��s��&��Iux��RV��.�1�+ز{`p/DP��<|1� �RT�qص���T1��a�	>%��ډD�]�� �*�����m��q�ĝ2i���O�Jv�qN�e<��f�6�ܓ�����b�bճ�&zrU����;�G�@��ب�b[H������옝����f��_j��Od��rP�)s�K�0u������y͓�w�����?�4�:RP���������>���&�W{����.>7'��=��݊��J���%{�7�UhzH�� �B�#�WP̽�
�#�D:�N���z��{����г�}�b^K�b�$7מ��	I��ڣ���c������yx~����k1W,�H����t/��z}C��*
��yPm��n�k��FrZ�҆��� ���v����R�ȇi���f�فN`�=v���e�.o'��*��Y����wt; G',��v�ӌ4Ș�+	TI�8��T���Д�p�Y_:߽.��*u�7e��h�)(,p�9�)��K�i�>4�#
�x��b+餎��oE�A2H`C��+	�¾�	�C�{�3�P�ڴ>$�y ��V['F���-^.��1L�t�����W�+�Xl��	_a��k.T@S*y$@�,ڃ.��p5u�L�8�qlN�q@�(�`����j�:�r�S�Iv�F���P ���@�&
�D3�g׺�iIoQ���b�B�F�I�b���&G�|+T�b8��T	La�J��������c%�*	��M�=�IsL�,_�A' ����y^���G�7�/L�� �Z�%����nd5���4Dm����٤s%e���k��)��q_��~�Q �X:"�M�ǭN�qH�F�:;�,&'�
��^|��\�2%��[�PІ��r�5�oBC3�|�{�9Ȱ/ʲ�!y<��c�o�|4>��ըQ�"���"���k�+�5%6ڌ��f�6AC��%��:.�g�@n�9�C���3��_깷g<4ǧ���O�q��-0<��D*i;�Ʒ�3�.��î������U���,��F�b��U>�f? 
җ��~)φ��Ѹk�_à�^�
�1���s�jh�v\4�
<��n���U���+c���4���
�����	.���ڽ�W)��1��6�
�S�_��P�´��������ha��ݯ��ŏW����ې��$7
�ɍ�������]Y��,h�"�Wt�WќN-�Qf�;݀œQ�]pU�>~n�oA�[�GrC�Mz\{j�j|]��M�)��j�������>�;�V�>	�ų�7#��E܉wƫsf��WJ����w�i�V��|Υ}}�<��0YP�S/T-{�����u��B,��k�b���th��7|��oB���ջ�e`
<�f� �@Ġ{�f�HI�
8��j�(�"�v�3Eht��_I���yw&�+���;x��&��G�\�u��{��s�.�K]m���	Z09��2�3��Z������6X�`�/H�ܴ�ޗ㤣��ò��eu��&�1��V�ڴ]���;�	�u��4�`��2:�P\���-*N��F�����ybi�#9EQH�B�z�3i�羐 ���X�Ś:wY$,�iti��p\k���0�
a}�6-<ÞGF�θ1�_�L�e{�l_&T��I6�%�hJ��C�1��JRx���x˝�`���H�Ri��@����t�������F��l��C!З��"��	O`�ʊ���К`{ת%+?�&������Ɔ�:����Qj�&[�}�V��7QU�n�I먠hE�����)I�;��+#�8]"Z��1���[�I�)X�4N`�����4��C�l�N��e׌�[�7C���r�If �uNXev��X$9�B��5 �a�B���gp=�ƴ�E��C[}��������z���)P�Z��Zm���܋��n4k��|������	V�; �a[ȆI}��:�݃�MO����P뮃m�?�m=��>.���Y�4\'l���D�P��F�c�k��Ԩ+n�_;.:�r��m�5m��C���D��c�ֳȣ�j�n�����\�)����Qk2X�P8��1r�������޶F|�x����r�7�tpV�)�p<	̈0`�Ίӈ��X�,�<a� 4r�
�L�+擵'�"I?���B�\��j̫��,��g�!Ib�^����J��U����f_TyTl�����Mr�π��Q�W�rm���uP���!�H��jL#������E�TWN�N�1KR�K[�tƎ;_�a�лO�����qD%��Fb`�����������XIũm
��Ϭ���=5S�W�o�L=ӫ��~�lp�5/��O�'5f5̰������i��8-�LU*GOb];����}UޓHH�\�%���,���ϳq�09���:Y3V�D��H�)�g���2c���;ݐg���2�y���ێ�&���*�x����DN��r7DZ���T %��{�[}^r���~����b z�A���O���C*D�ю���@��f�g����A.�e�$l�m��f��Ø�� 3��
���e�I���P �DL�$�7!#�u�ZEϾ�XU�1z���&��a��tJb��ᴻ@#_Y}\BTV�n�1T]K�|5Ӎ�;э|�y�3]*ֱ^7{Ia������~��.�S�=��	�۵���`����	�����~�n�	�ԙ�Or;j;�0}kς�u�&U���C@�G�ɪJ�w�B��NS�\@�]j1t��K�xB�Kj���y<�x�>�F�j�ʸ��d�=5�a��\�!-6d_^z1�L<�!)���cF������]:-���K�Gymw(Z��_@"�%q����0a��X�G�o�$5+�ç�&��Bkď}��r�)����������TYڕ��G��a21Yn�N<�ܰ�q�����������։j��$gf�G2��B|=�s/s�`<������[a�t@^8s>j�0sl8�u�O�.����]�զh��y	����*�I���Q �{X�M�t-~�̣P�N��P':�$k8�m�'t�aܣq��m$��N�14��h��!xE-s���k�۩�]Fm$Z>�ɠ������fm��Sa�	,���J�۳}�3��l��P�E�]e��O�|�|n��)�T
��>8�{4�gD��Q�˵ƲI[�L����H��Z���u�ǉOe1��~��l�XVK�<�nvCG-�)O3�HV�H|B�xZ�N}�6�ӵ�V�;g?�Ζ=h���C��%�I��(�27�-A���?��'WA|�:��k�2u;T;D��P�����e��Lk*l�%D�n�����;��(Q�T����+�w���1nQ�p��(��{�EMr9[��2Mɰ�p�u���@�hht�f!��g(��G{l�(b�(,J�.����RɆHϝJϗ�!���!�R5:qco��?�
�A��M����}W�B{��O�!�3,=D�R���^9pE;����6:�R>��G�8��%?��00�)��(��T����mJ�&>�1����ϣ�����Q� %)L��g{��V{���sjp^�˧�l����t4���Mx�=x��f����<X�5�dǕ�h���Q��m��W�!!���=�>����X��l��ໄ�NC�V��z���P՜�[IX��ɼb��z� �P�X�����3���Оe砮	�9>99)[����-g�k��7��qY1�;�X��4+2W]
�c�Y(��6xʷ�I��;@��}���^'��7�A�%X|��
�t��o�ȹup9�)R�6m�''����g����%�W�@<k���]�E�S��ۿU55���
�<V��[�d���t���E�C�kRUK���->��;aǷԎ��pJ��;up��Je>S�왠Mbn�rOnW%��g�q�� ����o�u���h�2Z��I���e������x�,�p��N����ߍ@�R߀�6�bR�p5����`�F<i�:-�E�F��1t�u�j���K�Y��Lr1�����C&��9�>|@
5��B>/a��6@�����a����O��rr�8gP�=:����}[s�ǋ��[����H"�B��D�}�7φ�"�	��E�l�����Zi`y%�z��Hz��Z���n��xi$0����TH���a
�2�u�_IEƌ���}��Z�^#�܂�P�»`�\k��V�����b�[ng~����J�Ҧ�K��md�i'��÷������]��¼L?{��0�^�:m�M����n�N��6��ǆ�]��U��*�z<�$���h~��?� �3h������3��IJ{�r�gUW����w4���5�z�$�T��.���S(qκ�f��z�o�&y��f�����Փ	�9��;h[��9�g�S�r�mȗ���6�3�J؅���]�))'>wX�!�$�r��9����ʺA�^�|<��>�Z�|�e��u+�X�6�tcz�/Θ�A�jA�0�f1{Ϡ� 9-D�B5�~|����e!�M�M0n`�p���q��6�!97yNt�M13�I�2�5t�R�	ؖ^����AP���[�y)*������B�-0�����'������E:�/���v��[�Ĝ�aO$;YD˦��[n4���
�ԌF����C�6n�F�,t8n�i�P�,�~`-V�T9f�m�����n���CC3A����
���K`��!������!��E���s���G��m,N�������1�d���$CI��� u�Q��GW8�YƗAT�*��k���vǳ���6��b���6����?ޙ��_:���tW0A�~4�4HX������v��^p�aM.Ϙ��JG6�h&��7P�X� iN.�F�N=J���i�>Vv�>jZ�eӮ�eeׯFf�{Z1����-�`��*���==���`ߖ��Oh� ������`�)f����
�g&wK��=��c � 7��'��{���wʤt�ֱ��]`l�V�e�N�@I��:�rQ�>���v5��,���Q�
�Q�R�t�LM�0s�����G�-HA���=��h�Lp������/�����	j���p%��2%���-O���79^�\�N�ê1�[�S	6[�~*.E���Q����$0}Ux-�2�ȕ�0�Z��扲l&utgSZ�i�@D6uۑV7�f�M)�zLa�ÿٌ΋�#� ��~ѣ1(v�Z��E'r|��[4��V�&\��>'.H�Ob*�+����a�6#￼0O>��Ʌ�p�	�3&�,8�[n4¯�4��l|)���Co�a���5�5.Dc�c�����^��]}ۛ6U~pŹ���W6|[汅U%���W͔F��಄�[~g"0ҽ�J���_z.َ�o�`=�H��gMଡ଼Q
$TӔE-8���kV�թ�I0g�?�4p�z�e�|���B�zTr��N!�fK-�E��NYƃ�(�H�9Ќws`��/JJ^�ZP]�@)ڄ��]�Oi��~s�h�q�Z(�����?f�M�ȿė�����0���h��\p�;}�F�1E��Z-)/4����-̷n�HGIm�C��C��hfW�Ĥ�@#���#�MFL3,��+�"���7�W߬�y`_��$t|#1�yَ1n����|�Ny��N�2ͪ�і��F\�_�q��\�);����2�m�ES��5�Ob:��`�jY�Z-׳<g�7_�o�Q����P�v�;{��l��Ls�ؠ�s�[{��V;�p�t��`U�����/�(�X������c�bK}� \ϴ!��;*TS=�lwU��NR�s��Eԡ����RH�D��E�RVؤ�6WB��w����4	�p�����!�@c��S3H�u��j�	�[�G'�">������?�2哲T�+��Z�"�	�y	`��}J����ڡ�}�TIԭ����`|,h������ņO&��VA9�&�2�w&ɩoc>>͜�A���ȷ�ϸ߸"��\���� 1lwJ 2�5sV�(��'z�F�<��(,�7�I-D��ڞ.ȷ��ԣz&>�i�%P�2�r0�9����~�< qlj%�L�i܋����g���2�_��EH9|�bY��gy'_b�/����k�52���
�W8y�KS#i�HSB �ͬVp<N��ڔ�I����'�11�NugN��#��#������Z��f8~�txB����ʖPt�vu�J��g�N��w�`�hNX�*?`x7��cx!M���W؆��v9:k�]΂ l���]P����1��s�8m��_�}��k�-��S�����\��f�fy�_��'\Nԥ픲��H�ޖ���!�w���Ua��N��BO���B����Y��Ma�l.�03fXx���jW@�a|�M�T��g<%HU��V>��p���m��$��)�8��xx��3���::Sm&�H��u�s2��DT� ��{��R�nS�Ly=��6�C��L��9٨�B���ԑ�}�6v�!��8�ȯ)�Zi�
ǿ)���Gh{֧��u�~�J(�}��r���:v'X�'C(,��!! ��_�l������>���yUj���"]�V}��i�
P�Gx� s�mT��U�I�o��������">�� 6*X�����2Mr��;V�īՅ�~ ��A}A� nO+&�$��am������)&��9�pڔ�(�m��E���U�#�S����TI��י����m��Gh�C���De�����y�T���9{a=�f�@Dڭq&rR1�`�{R�V�<����{)1c�^��L��?!D��P�ǘ���1]K[�U�t���k�Uȅ�3��־m|U��c<
K!CqhS��a�w�gqK��p5��Fzk�P��� ����J_�}�A=�_��[�����.�<r��ۢN<�f��0ⶹ�:�i�	dQO{/����t�,�+Ä��K�7X�q��c�~��m�5�$|z�p�$t�]�g�7�1�C�%P���7���i��+��p��ֳi;�af�e=�N���%������cnV��֗Z��j��+En����`J��EN�\�@?��߼V�ңL1J�*e�~�����"J3���*��G�J�OR�ծw2�D�pK����CUi����������$���]����u���<���GT�i����i	��_r�۪ϙg��̄��	Q_��2,��P� �ll��L��h�H\�]�ً��'�ԑ:��E ��YF�)�mg#�{qOZ�.!�$�mR��=ra�f��Q%�rzu�� �d%�F�Asd�=�?]p�cCZ�c`٢t03wpGaM�֦{]��6V�0/��	�LYh��Y��	-L��W�^�K�$���c�����n�Dțk��_�D�'A?�9
��7��Z�����0.4
F\��Յ�j�t�V<��κ�V��	).MW��6�ָ���q�F�X����+���n�|�f���	�9���$`�j��>��]@��x�[+\�Pl�yX0�rc�����@).a WV{�| �p?�^�Tm��% �wCRϧp������-����),����. �Jh�C�Ǯe\�T�^d�J=�)�+)SBcH���� ��;ƶ���eFP���}E.?4K��-x�,�-�$��Ӝ�]�c.I�7�h��{ �p]E�|k�z3^d	Y���8$��G��+߭�(���=�+��,�C���j��'Krwj��K��9m%<SZ\�
���"��@��ʄ���׫�VI�m�P���ZE;���s����yS�0%�6�.��c�tC+0�ؠJ'�?I٤��ύO�`M@O�j�}3�0;}�z%K��ՠE2�n��u$���C�:~`s�i�	�<3��K �m�w7+���J���K-�gէ��ɿ���Ri̏|r��H9���FG���|3�Nf9�M����w—F���YX��-�{ϝ��+� 2���9)���/.F8@����mF_�1�R�����{��*�3A Be�\�~K���l ���o�S��ƿT�j!�,U#O>�6����d>��	}ÈF�H�<�M����6��ˏ�]0vE��y]�?���Equ��S"���(����I�G�u7�烵�;v��9�ɻa��i�P2>��}"��wz征>0�إ���vx�kg7�o`�X;��bX�Ku������9�3���9a���E�6V� ���$p��Q0D��g0�L�̺�	�Rć� ������t�_AB�X�So$��\2)B�8�����͝?���"����:��61�J�Te�h�S�fս�f���ev��Z�iI]P7^=+1��K�*kx�'��Hkw�g�+|Gg.%�����q��T���pOu?��_��\ڨMG9����gM�0�d�?w�<H;-���M���<�]ΰZ�<m���%7��]Q�_{�P��e��Kֈ�;������C��JI4��E�!1u/�z���H6זz��@�"ɗ����g����+��WG��7��)b����K�K���9̄��CZ¹T�pf������4��F����"xY)D	�Ԫ��CXvM�Q���q��i�ޑ�/�x�	 Z�^����R^J�I��)��h��o�3��Z���P�w��&�-%���}�A�Ҽ�C������lOdw�O>�H1�bc4i�A�arsc����}?r:�PnفU���?�{j�)���S��;��c��7	�3Gi��� ~x6�vSom�)iW��0N��4�HSQ�#�� ��M
�hF�j�2��EOY�u!��X�DȎ&�hVb���r]tX�ZX=�'%�"�6x�Es*�pjr݇mׯ��>p>���!�=oю$]K\\�ro?j�+�^DUZ޵c�/�	�J��a:� rHP�?42�'y㆟�)��U)����Ct	��:��~����f�A*{G3f���ܲ�!��{�t��T�}�4j�������-��[7��L�7&�͠o���,�����H�Wi\TX�&,N�B1\8���#�x�zQ�l1z���J�Ԧm�i�->�UnJp�N���B}��Y�i�=�#-��:��5˼�ϵ��4�`�uC�4�+'��G^�?Z��j������3x�B:bʲ���H&�P�k���y�R>�S��^�3M�1��8��{���ri��/��wM����<�e��1���W��&�vÐ����v	T���ԗ:�B�	��4&��\����{K�:�\����"\?�\��Fڟ$��u���-�ҭ�B|�tKk��8�5�`n)aI�C��g@�nƻ�z�o�@7��{و/����j`�N唲!xM3Kx@�%�n��ɛ*b\kL�����0��g���R�����I>����x�4J���[�� n�w��R'����hϥ��li'���V���2��^b�9�?��󚻱��߼��_�0�Ju�[(i��uH�A6��PsV�]g�،}y�|U�[�m�}"����W�Z��?��b�X!�V�B���y( �*oݲ�T�#�r�,cp_���-`��]����Hy��QbG�>t�!�ý�6���@�jMF:.(�+l�ז��X.{��W�� �EN@6䎚��(	�F�@	��:��7��1̮�{�Qzڎ�^�5�!	qI��:��Xb���)�z�^�hE bn�F�����֬�!�xk@��֔+j��P㟄۵�w�V��P��S�T�9p�aG�74r�����e˭g�E�~������
�u�����d�Df��fqc����,�mdߛ���ؼ��U�<	)������51l]����Jdz�U5h�3��xK�ވk���_:CM��iu�8ŨsB����q�S�|S��P���?y���ow�ug� gK*ͤO�9��3������)���ye�\��m�k���O������A�����@�����q�D�_�yBW=�B\���K���.�A��Z��y��ڍ����ܷ���0��Q�u*e\�[{�Hu?����z�Ij~�t<c#�bYb�|���ݿ�~f� ��7ʜ?��u��A��F�q����+��t�������`w���|����P:Lk]�p`��ګ�H������T=.A@�ITI�F)�)��.�iF72�C� �qAi�L�s� ��d���>k޺%
���+&E�������8	�"ƊH$�L\7�vGl�$ `��x��z���J�D׌��p|@W��,�\'��/��G�qSl�k�9����Nec��u(z����6�����2���W���&CX�jh�/L��[kXI�#��E�-`�Y:7�cx+a�-��4�L�A�.:�4��@��U,�'j���˼+_�`���lV�b�o[i[D�`����W/3GYA��{�L�\�]i�q�����笙�N�Bx,�{��DD�L��O	��C'�ֽ?���+�)�KG�s(�׭�; ����p*�h8m�Zm*�@�.i�Bvn}����>]�+9��m�U|O)/n7h{�R�FPN��V�$��pn�����C(,�����8~9��o��K�V���XK��<�7i9)�_L"؂&ۂ�"���-��@�xF�n����z�/�G�|�Ż��:��p�H+h�O�9���V�v�*?�R}��N0��.q�Jp��܆�Dn��x귍�al����X��{����x�Q�/Z���yV|�B'�ԭ
��?�H���ҵ�u� a�6���WX��h��	/�Av�"��Y0iH���P�Xv7��"{??z�4FQ?[o
��zؤ�IE�!�&e}���=��x��4���+�ɠ��>:)�F��?��[o,��̇E����H ��7b���V;�(�V4�~�~~|џ��ٳ�o9zn����j�kpfP�ލ��HoS;CT�os�G��Z���������J�A[��tiY��%���G�6B��a� i��ook\BGߩ*vh5F���Ȓ;��7H������$y��M��aR��R�5��I�@V-�����}/\�F�K���Ǥ�#1t2^�VȌ� �2�jy��S%I^���k���qhF�!$
�yJ&�R���0��ge�Ah[��@T@��@_q�[ D��79�j̨�q��`.��P<�'S�����r e��@4>I�M�y���M��8K~�o'@n���å���Q*Ӣp���P��h��Mm欼��� � ���n :7`f�&��}�L�Y
]�N���g�>�)9�TgE��<tK�\�<J�+�l���_^K��B��lt�KܘT�Hjnb�=,��`>���N�;�ɺ�fU*���dE�er� ����{�X��H?I�Ԛ5�u ��R��-���a��P��O�6���>�&,�>�_��d�+��3�E�W8tTwQ1�槸c�Ibލ�Ҵߛ"�|Ǯ!6t99C�{,iB%��uJ�^Ժ3�D}�t71��t�eE�]a�iV��[KJ���s�|1}F#x�Oa]�aϩ�ɭ�>��6�鉱���G�ǅ�b#Ϊ��"*-���R�I�j����PD.�r���}/�P����>���IEȱDI�ɕ�����ڹ=o�3�^`����{�`����/�/�פf�;�~��6��F�u@��YL��+Ht�{g݌L"Z��
�Lm9fפ�9Wd �h}ugA�e�˾B(���j���vfzE�2�:5��پ��\A����!HO�4��2�����]��$՘MY�L)Ս6=S|\��c��_:0��[�zv�ؿ9���k�Q�5� qN2�	��&����H����:���n��EF�]����6�N���6��+��ޟɆ�
�k���NFL� �)Bϕ�C�GL=��{�da����ã�pM!@�꿛;p�`�Yɰe	�"3,�� @���p2C�M�)���p��=�&�����΁��b�q�Pl6���&k�C����[��d���.��խ���ʗ�)q�����Q�䦄�k���D��ǮDtEgM���U�.�L����%<�]H�m�m<ǡO�~�Z����>�3�&�8_ya8��3Į �u%	�.�L�����nH`��e��/6!��T��<��΃_]�L*��Ү��-0l������?;����xmַG&p�Y����螷��l�k�T�|����o/���GC�2���8�N�/��d$X��L���,@r�ܲ+}>f�p���4�����"���mЎ5�c��]U	n�j���"�ZE��P����ۆNt�T0	VS�JA'%��U�rN[^�H��p��}L�? ����%��cJhO�x�����Sэ&o�=I��Ud�r�Hп��&�`:���y3G|�AJf7�H��W±Ȼӈ�f�F>o_��HW��&����Wo�r��퍺�R����YS�(I���bt�J�r����L�]x�PŨ;��c0Dj�4Ǖ��8�p��O��`�E���Î�W�DB�����2iB�O�˚���#����p�T�{�=�Y��j�*qo>G�8�����~�x�-��G���G^�ׄ/����}ۄS;(�|���lvg�b�hv������r�x�����Te%����+i��5+�Ȍ���L!�:�T�XZ�r��2"ף��-����A{��EB�I~�3���#/��y^�FC�X'k˿� �y:��;	b�C�s��x�.E9h.?2% �;∮K)�B7��C%y��m�I��K��om1m����#U8*�f�����;9�.��ci�i�4�W�C�Dԓ�[�vJ�Oͩ���-؄��شyj3�3���	8��P��7��ѱ���`�b%���6�8[1���[�W;��	̊/�Z�Y@�]�Nj��%�pA���`��Ćg��gv�𑢳Ce��z
�(�|�K�A@�s���+��0��!w�u
�Ŗ7��;YAd�u�āc����������F4��9J��$��m����
ܮ�����	<a����6��F�S��L���\w�w�\<Z�Wk~�ƒP�L1�!4��B�wq�a�%�p]x3� I^R�8�iX�r�zˌ3TbB��f�%�Ȕ�?�]��a~޾,%��WVH)���i�;��45�ϒ�SnN���t�x��։�֑��b��.6ɕ:�OD�pk)��l1�/աt����Kƒ0[�޼�;��~�c�\���x�$p	j�un�)A�E��JpRM��0�}�v/�R$��n4T�Q@�����+W���S$Re��';r�ӣT�65��8�=�1� {�2�÷Pg����q3&�4���P��B��Y�i7<9W��@���h���vH���R��&Uw��D�)�J���=�F��Qc6X������M�{*N���ԩk)�;*����Fh`���dJ��hM���E�J��X��D�v;��.�
yo�.�Շ#���nj\���'�=�#췎�9\�A&���cE������a5�+5-��D�I�7KK:�yehA��C��֭��t���4����3Y9��>t��@�w�|��
����Kn{��5H��ģ	�oc�	U'��-OMj�G��o4jp
Q;�f>�R�ӫĽ�$W��a���(��
k�� ���f���FӥÜ����ec��Cs��̛,C��w-y)Z�dݧ��.lj9(��M�8�J\����/ضɠ�ӮvrѳKЀ�L~/�����&�	P�F�"y�_7s-�=x��`{xC
�*]2S�Nq���e+]Ο���O�K���/;���M ]>'(cjZ��p����
��A�t(�d<^8�
��c�p���O�{��u|����-I �_��ɜ��v�	,�ʜ5j�'���F���0�BߌV�w��� �I�P�}�N�"�DA�f�42�i���7��»H�@�GJ+���ﹷf���/��=�+��W]D�����ɣ�YH���s��q�h��pp�'�H�DI��.}�������e��Iun�D�NySe��P��^�%ؼW�'�~J��X@�d61r^�;&�w�́V�<�6Y�O��L���RZMb��F�����Or�O �h���� k!ݕv/(����)��6��u�o6�Ύ���7��%���*�K��|xd�s�[D��%��ib�~^�s����pm����-۠�}��d>l�3=6�?X~Ji��R�s�'�
4��<*��¸�U1K�
�j��:��j��jLM�|���/nj�lį6z�	�-�	�xj�p>��^�q�ݢ��Kr51r��"�sqw�zBm��%ս"�:�f����8��0>?�^jN���Y��M�	�E���j��Xs-�Z��r��#
|��%!j�}���P�%:���3�R��;��߭��70�G@��������ޢp��Q��R�t�:U!d���V��4�(��2���
ζ��:������"+��y\'
ܤ�M9/�T���`?N!F�d=���A�ɿ�OQ�������N3���}mr�G�jVQ�Et
��/V�?�pm_��1|�{V��NEɣ��Q�:Ȣ��e�4�B��,��C�,R��Eo({JNd
� m>ɿԀd =<�+.�\�]�. �1�=K4A���l�<O5�u�4R1�����?�ֽ˧ �s��z�k���T��>��컃a�6o�g� ܖ�h��l���g�覕n�!��j�H���ޛNa������EQ�����j�{¹�R���ltJ��G.V~"7/�Pn�%vp8;�~�5��Ol�?�r|y�i�R����H������H������H��b5׵%�Y��]I�3�ѯu88�F������Z3�T�R�<Q$�0�af}H*uj*��8��RSIt&��&)	ŭڦ���3��!��ݾ���uY�B��}ME��C��!´v2.����ފ��o_B�ܦ���Ku�������K�9|���W9y;i�@�K)�Z�۫w����6�i�Y��?3_]/�8y�1�R�A�5��=�$��D�,�mZZ��v���_��Jx�=�j,_����"ya�<���t��<�MRՉv�pن_n%�`�$�d��rϩ�;����HaKO~�I�K����n��pc%q��c�䁶�����*nP�n�\�Ū>2���L�XI�e],H���d��Nd�ol������\�ⱟn�8���tҫ�X�n�+� �f���[�6K��V���ّ�e��>X��Rl�0�AՄCgAkjn��c	���,H�
~&�҇#����	�"��(���9�r��B#��'�ff�ibf�qb�U�}a��."�Q��_	�z�\�<q��;l��U�3�Xu��� QΣ?�3^?�J�,�����M�#�z�ȝSp�f����_�r)��g,�vQe�~�m���<6I�3SK����Ƞʋ"iZ���Y����.�����4��kF�N�iA���ܗ�����5��VA �`N@/d���۫�nS=��K�ݲ�9����? �ģ���������Q�E(H��&�=��A�)�(��;9�J!��L��6���P�I�~T�RV�Z`�c��Zm�9����i{o���2�D3^S�vC�~�p�� ��T�!3��:Bh�P��<Sq1	���邲�~X����?g�w�=�L�7
�����/W(y�ݣ�uڎ�S%��A+f5���L�ҁ��⫬*e]T!��%��ų�,�bC�,��&�?Oqf��}�����@�t4���Uq�4#�������Tя�?u���sknq8��S�ЀAm���~%��n�IҲ�q��X�e�؉�o������\�������8΃}	�h�z3/�D�<�ףV��/�D+�z��1�i�0�5pv����jY⎝�A�L_�6�bN���[o��J^�-�&~��E����nV�Q�f->9���`')ɹ�'��_���L�q(�E1�l���貰N�����={�E�Ggr��)0y��cL�̌ƀ����(��J��:ԥ��qJ���8��l�]��ʉi�f�'��\���*�x8���w��|^��e����b�W�,~v����dZ#靝�+|���b�[����9P� �:�ȉPq����A�\E���P,�+o�q6:�<WYg���Ǡ^���*�.�eP,���
�Gp����en�$t��j��j&ٝ �cV�J�%�}��w�ܼT�勜�P�hi��W�!�6c��a0Ͽp�C��^ ]�J���:A�nN�񒃹��y�OPݭ��ݣ�8��Ļ����(���W/�n�~u@)~n<�'OX_1H���幝��B)��O���ݶ}�D�=�5@6��G��6�k�,�B;f����PF�W���}�W��� ���pZ\�;��{ }�粼�������J���x��_��v*�O�'ְk+�m��/�}��	$	k���Nwz MA��k[u�(U-��$Ͻ�yc?�3���wˈǐ��P��%����d�7[��,�s�}����Mew�a��90�B`�??�z�Q��3$�ަVJ�����̖0�j��m�� �+%�A�����&��N�>2����*I�	��2�H��M��٘��~�	'椿SPy���=�,��_��D�N�%�%���?�u�Lq�]��o�J�꿺��̶h�Q��G�b�!M�h�W7y�JFi�n�H=�XM/�TN�̆����G�:{�:�b�'	�ݤ[�Ԫl
���%x{%�+WN(����ԢɅ�y@��s����f��iyX�>��<���N)�\V;sR����O-Х8�O �)Kٲ+G���O��对s���������Ƞd�Zv�8aEp��Mim�3+̥ϔ��#kzӒ�Wt9ë"�%�!���1/c�U��31h� �#V�)�H�]�oK�w�st�
�� 찼����g�_A#�w���� ʮ�LIV
R���/��>�Ou�b@�KF5���,�$��;�����+^�0�8}��'C=��LKM�<��U��%�B�Hx�P�ۀ��I{�>��-��89;��)�}�-��D�zf�9:��D�
sHʁ�(�?)� ��s�Z?�4����vw�7� w3S5ǁ��0����ٱ�'t?o�Yn�.݋\f'�s����X�n��I�츺����}�J޾q�ձ�T�)1/�H��l��@��z��L�v���NZ��!�c�Q�&:=�I��(m�ew73�0�4l����`��%R��R�����C��9��0�Xx+�/mz�f�I��]�ܡn�x�%�R�B�}`����]]!�X:�FH<a��=�y��lHL��':<n�;��u���l+� �2�TT��k�)ۅ�#�1�m��)
�T��^�$.z�I ~w
�S���Q]"SI�^n5׿�ڹ��Α�ZG���\��>�*���nn�m|N�1��z�J��a �~���^�)e?�c��F8����5�%S`���2�،�ĩ�S�H7��<E�Cx;�\�[`Z���z�|J|a���ՙII�G���Y�&��K@�o��į���e`��$ܳ��NZ����"x�Qlh;��e�YhTL�q����Y�~O�D��ߎ�>�����T�{��@�u�'	�',�h��l^zt%�D!�S�$�Θ���j����S�,���
�^�Ŝۥ���IU?�Զ�����%��8�\��ߞ"5�Z��6�]�g���*7�$Q�aA������.i]�"c��\���{�Î^�!�?���nJ��3l���|3�^��Fm%5�Y��%=�^�!�n\�ʾc[�ȧ�-o�Zn%�k���j��q��u��/^d|/����~e�wít�W�j�~8O��T���+?g�ܿ�b:��1�&�H�n�;��wV��~'�X77򁓡�r���7�2n!�4�ߍћ� _��c�2�v�����X�����nN9z����ڌ?����^]n�W�1����y.����a���0P�M�vW���Z�]�5����SP���`(S-6Kg����-':�L��4'g�q`0�P��a-��H�����?
?� .��J^��� &f���w�ڇ��[��	m�U�c/Y{�e)���L��2�a�}`"5&�*�8/	"�)��L�0f-f�z�K���l�D+�l����JS���V����dU���d%n��J�V���=s$˩�\�(��397�;(8����Z$n:j�HG�UP1�I�HF�NऐFȭ$���\�Nd�@h��}�\d��w�E�&�#������?~�-�q�?���/at܌�5��`���z��F¤Aɛ<�g��@��5�vy'@��8L�Y�o�J��&A-���-���\:�����g�P��Fd�(��j@z,K���#;��Oq�r}�B ���t�ի.SK>�y��
!�6����J_��qqhѼt�UT�.�G��!Za����H�.7��F�>o�<y�o_	eǧs��c��l���,4�Z��!��;�3�<#���zx�����?R�sr�9y����h����q�s��	9�Í�� �fd�8�8���xꜙ��2�|ZQȬ��Q�+n����:��Y�5�F�?~��w�a�����F���<3�:�?�E	B���W:,��(<j%�2��s��ٛ������u4a_�C�·�X�`�ȏFe_�%6���=er)�of|�R�qz%�z,��24s���!H���[�Ia����ă�%K�zp�Lix480�6rR+%�Ź�cBL_���<L�0�*�:�!���)ۭ:�iQ���/�fЖ�&�+?�������Uc݂nL7p!�7:�MvC�"cwZ��q��Q@}�+��X�AO������g�5�3/���No���I���$5��3���g�`&]�I��[���t�4�)�B牪n�q��!�	�2(,���S�Va����+��'S��r��T�|��Z��33�N��&IN+��8�Umz7}�6��HC^M�&t[�e��ۮ�/B#lt�(���Ir�e��'&�<|-�L���
z�6��Ց�iw-6�!����E������MJ��I���8D���N��f<:�������cQb�K���i�#�H�9��+B{)�ZV�G�%��Y�F*���Z�6.�I�um�y�P6`Y�mYJ���Z������A�I��i1�Br��U�φ��3K,@��	��%��A�@dQ����}��T�W	��~ǵBÖ�שׁL�2x<����#�̧g��>!���a��l��L$D!f����#���y�ћF��'�><����%�Q,���k��F���w�C;��q�($�t¯���5��y֐�:2��>��J�nT}��]m�c�M=9
d"�ֳ7G>�w�5=ׅ_�-c��΀k9�n��x`e��!`�"��q{(X�8I.�Z�W:9`��������r���E�I�	�|�zU�t;�)ζ&���&rk�
���G�Ԯ�wM���~�@
��!�����1f�z:\Dt5���j����3���̆�������co����̃�`F���/k���Vr^�Nת�@�SX��7��ax=̓����+�E�k�?�����N�����\���u x�B�+񀹓ӫ�X!KS��>9r�����?�;.��e9�Z�9�[6=	�O8�!=����	��������+=�J�u`���?���c=�?����㱚u����WA� �Y(P=���v��Th#�0m��JZ*TO���Q�l�?��~'�#*���y��D���!-�E)ފb�>.�;O>$1�uz��ڢ'_�lF�2���!�;�����eO��^2Z�	:��U�|}ity1*�P1���?u�H�Cگ����=�z�6|��b�q�v��{)����h:�kF�Ж?b�T��*�������-d�&��.�2�;�{�2<H��Ct F%�������5�.����YN���G�b��G�#�?��.-�5�o�yd�M��
�q65.��� �/IogDF��4ຊ�[!��b<�����@��CN�c��/S���>��;Q��I�1�{�ӌ0YT�d��ݛ�)La���ֹ�zh���f:I�∳�Q�Y�HQ��/C��n��D�Ca?<�i��ڬu��6H����'�o�gn��Omڱb)�j!Q�� ��,�b#w� �o	5R#��v�ֽHzm|P�W=�x6^��ص>b�s������Ix�Y)vl= �!(��6a��ȅ5˧D�Dpc�@&]A@�d���"@�i<Y��ō��G��|�X',@QÅ�Ƶ8�9�t�?(cw�Fp8���z	a!���Z��2���l��x���ܾD�
�_�竑��O��E3��6�+�sFD���`��xX3QҿDp���҇��1.ہ��ф����u��bR�#;we��ќ&�q@��/�MO�XT� XZ���%E:5B�#r$_N?��爝��p9ͨ��4��/=6H���CFK�~���������oG��؁
���7��^�/��DI@��_eϥ����x�<O�t.��큱_d�E��U�\����9,�в�2�9�~u+W;�m/}��K��^�@��w�l����I=�MZ���!�b�͸%�Cu�ɘ��"��潣�՗�ŗqJ�9zMW/5�7P��Q���5 o�O�eF�R��O��m�����@~{֚V~۳\��	��Ś/��Q�n��8�zҫt|�*9{N�%o@���)����P�6��Y������6�\~��ۭ">=�e�M0�Ү=Nc����,��^�`���;Ա������J�4��С���������Y�wʺz;���_����?F����q�ͧŞ���E�vv�2�>����d��b��!w���M i�{^���%� ݜ�`t���_�Q��B���F�����;�\�M�JD!_2�!Ŏ��U��a���m�\��q�-�	��ϊcVo�R�;AG����(b�A2�Gs�����x��,R#�F;�\`�.t���+���i��p�*`�G�|������sd��s1|Ea�d�ʩ��s7o����[!��xk�v¦;�ES
��4�r���b��-*�� �)�eϷB��X}��e�*V��χ��`�����[.��P'n+U�1H��ذ���ԇ:��b�������P�o��=����rm���$�N�:�`ǂ����~j>�KbY��D� 1�\4g�����K�m�	�osAjA�,�#�N�r>��9�_�*f9�u��7X6�+�(��
W�8Ѝi �D �����Q`*�)]�޶�v�V���,�#�=���Z�^}�Y�U]�7⡉�[*BD�ٮV�:���h(��)�-�	P�[����`���/�T�W>��j��v��b(�.���	GXx���J�Lo�J�v���n�Jϡ��#S�'���Y�Q��5�)��{P��ʷ�a<+�H�qR����x�\��P^�Dv�q���5Rk+|��Р��i^;��g����K��n˶h�Y���c�;�t��E�~*�q�yK�	�ǒ��-(̘u%��	�7g�ȅ��>/v7%�������2��Z9b��1*NK�Co�E�e��U����@�^@Q����\i��e*N� !�q��	��-�8�@!`���M�d�>b}�
>``:U[1!�ӗ�����To����ܞ��wGy�~�����B���0�}V��^I��e��'�׾j�Mj���s�ß�?���<&5��$f[���@�Ws���/�u�0�7��/�	��?mƻ���6$�w/+�0w��	S�2Y����T�9k��n�v��^o�_ee}�^�|�����gaDblӯ�%?;g�����.�"��yL�I���\@�~�|]g� R;H���^�)N�.�I	z�Z}aj��X��&,#�ne�9��N���F���_3c�q��;������~�	�����T ]��e����
�J�U�4Z6͗���h��wɋ�y���hsڽ��3R�0��u��))?�{���o��Dw�6�W���
�e���j�tք�7!a��?�5����v<=����K��~;W���.%H�;�ՕڳGp��/K���k�P�(]	|7��(�H����~��h	[:s\:��`}�'�
�6io���U����-\�(�����k���N�*&�E�켞 �k���
�x��v�i�����;�sy�ʿ�w=����#r�Y�O�Q� ���@n���{����}9�! ݬ�	�0v�R4�|"f�9|o��?�,��Z�v{���AT��s�Ki2��TW5R�CcU�:����#��B&Y�h%�%�_,�Pt��|�j���KɃ�5�e,3����/���
�i����\��ed�\~N����X����SiCd��z�xV&�_X��@�S��uQX�!�����)�>	�̉�n
�<�7	maB6�c�?�(t��r�čQϖ�9��4r��߼|��f��3���-6
�R���}���em2�9�����..�а(=X��>��4]Q@ւ����[YN�SaK*��y����bm܀y	��~:ho����E��%���'ę�Kt��R-�%�%&� �Q����6 ���~�Z_ͮ(��B���'����������G"U�+���6{Ľ`�� �;5����N�����˵6m�p�?i���Fn#
�j�)�"b>Qz�K�G���j�&�·<��2e�Ї�'w7f>�WI��΂{�,�xa��%T����@��\�~�)!�|܍����b���^�~�wpc�*��t���7����J��S�I���� ��"��f�s��Q0�\�e�$�0�ΘK��5sX�Ω�;��{<��?̫^�0�G�B�[B2�	OB��"���_>���셛r�+����߀.��_s�fٱ;E��1qu�T)�r�	36�)$-�,C1�z�s�=6�k�R��ɩ{���U���d(PS��\k�^�TP�/��@l�'��c��>/xd��?U.�N�r��D)1�~�Ty[qL�T�R�� 9�H��`����̮4��t_����k1��	Q5�Y��GI/d��vy ,�`C��ѣ^f���O��Z�m�L%��,��!$[|S.x"XĪ� b�ӛ��l�����JY2ӧ6��cTV�#���Q�4k����/�~$>�13����g�h¬P#�)�!��5�3P��q��S(����[yr�5�7��ufȵ�L�c�7��i-�D��I�k3�'Y�\�dI���_{G$���)���A�x:C+�}J�r0сz4yx�Yg&���/MBF&�x �sO��s���鮢y�LƤ�lbqX��2H�M��M��3l��+%���}[LY�(]�=�}L��H�m'�ǹLHp��f����˷����]�q�:L﮷0�-�����#b��;�,�N��GӦ.on�n-g)��|�Kk��KX�]�浓�&w���ОS�強l��F�׷W&�@]V�Zð 0 ���eɑ�W�o/��ѹ(�5-�@��ޯ"�*�xÎ eٟ���:��\�����sG�A��C���ֻ��S�?����C������䃈g���/yYG:޼R�����k����̇@kL|�G���Kژ�g5�%���`K��;Q�ҹ��V������Ӭ�]∈��c���7�a���ƕ!���σѢ�t4yi�g��@�:���ͽc4Z4��ܥ��<<�0��D���Ʌ�5��9ֆ�0����kTt� 8�g��L��E)�J;��l*�Xr�~����nN�c�Y��M������i,���<Q:41QDE��J
�{`��ԋ,��ċ1EX[p���킃�E�*�M�U�W���2����g� �;?��`�,�K|�*�<Cp����'��"�7B�$�䢏���p�[�'���J����V���kr�q�}�r10�lTd��|ň���n�:�=��>���2י��eP�������4�Ih�0�-��׮��r��@�:�4z=jhr�ZV'	�7ߒ�3Cn! &u]Op��@w�+�V�Ɩ�9�l�C�B�{1슝u&�9{�� Dks����6%��n,���#0�Fd��}ŭ�'�����D�W<ּ���V������N�̀�]�֦#���:�L&�o��C@��~״'�>�<��T(8���~U�g�HL�|6�=��V��i�[�	��O/PO���8xwcY�������eDH�u"̯34q!�9��̰{��՝��:?.#E�I �X�fB�n䍰���.G>��D�� ����8v��Gs�'�$Qw�_� ������y�tj"SH�u����XF{�B�9��"C���U	KQ�={*�U��+�0��W�Jk����zXߣG�ӱ`�~���}�6�4�8æ\L
]�F!�$2��kD<�F���C��,�����K�P�A}�r�}�#u����5GU>?G";Fs��$�z�b���� b&Q��L��(
��%�Ϭ�htzŽ����5����խ?(b�p;<FWO���,�t���Dd������)� ���u(���?p[q�~C��5[[N�Ax��Si�횠�wj��s~�꼼����I$�ޝjq"]���2b��^��޶�I=�uuu�iU���a��l���ڛ����ڳa���Iۏ!��O�zRg�L���.ɱ����G.\�������xd�P�w:�`�(�XG��6{���> �MC�=]�S�?Ͱn�̽I̱�y:��1gA��>�	�4��=��NE4�²��2�1��Ƽ��_ǜc+6�f� r�SL���\ڙ=�<��-S�1�9��]2�[�#������2�׼� �> ��8�X֯�����ac�"���?�|mbC-���ͷGɉ�*�P��ߋ�Q�D�M���d�����~A穇�y���<��';	ȯ\V�������| ��)�� ����%���К��IwYH��^�WG�n�8��/��~��Y-4�̉ngWa����-�����f��j���	��Re�$�'<�<}��-��$�ٶVۉ���֊�7 o�-���u}�'t�_� ,^ւi'a��6������<�o/3����Q�NEp�����@�"����W��8H(X�T�,^6�贤�:S��4�S�\����7^%$�p����0�A���U��������,���� `8�����+J��Y�'���Db���dw7��sD�:�unyd��j\��Q���l?i$��*|y����
&��A��p�Կcu�<W�S���Rtu���iV��,�~oo�-�A�-d����e�O���^wߕY���}�&��ԕ"@���	[������Ԧݣ��i������Ʋ�9�`�`��轟'��>jz����r�W�[5�؋	\<��|�}�GԜt��Xz�3��6�$�6�����B��0����'�Ȼ��`�A�����~+J�my70u�,A�d��v�t�&h�.@��W��e@�?9�����p�ɰ=6�'�kt��=ȌS̎�0M==�n5���ϖ>���ў����~É�M�n�bp� ��$Х:1)�Q��t%����kd��~O�{�1�QQ�t���K9��3X�?!̇47Oo+"�����9��ywi�:ȯ��GY��.q&ݩ�����o�?8��Fy�Z�<���n�<���}��)����h�O
�w�{�]K�����C���q�Ag:�V��[NF�p<�e��%Eq��G�E��γ-�v�roe|�,�"�A�1K���ȣ���2��{��1G@<�{��L�`�%6��ħ�A՝��q�1���;{��r�W�ug�.��(
���~á%=��"�\�H���s?������_{��`� c. H`I�k)à����u�����b���<| �Wز<Ӂ����h_��rA׮�x�	Q�?�2�`����+�GK����y)�A�m�|l�7$������~2�Z�t!���'�\ӗ��8��Pw�����B�s��2�#ސm��;Y_f����:`?\n��ӟzSɅ�^a�!%�
�!{з�dDģ<�����g��hew_��@U:�ˎ����������W2�l�/z�&�>Y�T����!E���Y
t�6dݍ���s��\5bb�HMrK�5�Sx�脤�����E� Cv3^����串�d+���Y�J�A�ܟK�1g%�H1��D#b)�����ߵ�0
�^�n�+#r��.{�<�D0����S�\�$�)=���=7A��I��/5y簄��� w/ 
����~q��|���ͺ2��Gj`��Nc�R�GY(b9�n�׽V/1I���{R{4�šS(5,fMt����i�*���M����}�e�����m��	�ޞt�mo7*�==�#"u0�O�גf�.��d�:���Ɖj{��VuY���WKq�3�,-IK�]�q���d�q���11#�˶8�G^�'��:E��dĄ]�tq4��z��ݐ��d�{b�� F�x����D4`q4>l�>���MٖbX�t %vaF���͛^������m��%G�	�V-�'U;`������^1�;���@/�@݂���pz����[�V4���� ��	�;��#���G��H��F��M���-Id�P�.��:�4������-F�	��R��������g���pׄ倏׏0_Gj�s18mg�AY٫�ۛ<C���C?U�e�Ϳ�C�>����6G��"��b\�qLN���b�.��Pf���R݂0��3HY���ԦU�'W,���ye���:�B:k8�z����"�,�!����:��/ ,Z��p_��ӌ�i.���Ir'p�p���*��dn��@�li����яëz� D�9�?�P��8Y�"��.�%�MR����`
Paئ����\�p��mvNZZ9<X��ߜ�ce�Z�5����/�i����5��q��E��a�X��l���O��F�ed*���&�]����Ζ�n����<�E�P5�<��
��X�P$]����D�i������Ȓ���z �йw�L z&M<�-~�����,ǭ�I0�3 ө����I�����B�����e���j�
�U^�&����A5͔I8���pMK�k�w���U�~BAZ���[�#3�b�6"�NS�Hbv��7X�ABA��{\G�F�H��v�S�/p��2�:гz����R4�]ʨ�x�ı��'�MHh��s[�-���Fiw�ս�\�d��3%]̆;S#Su���̽�5��\����������r�~�S0w�(�.Rw��VO�h�oF#J`�Z�	�Ӓ�XnzTE�U
���% �t� mJr`��\oR����w�As�t�Ak��Ā�w2:�;žs3�Y��~S�A���n����l��2ߌ�d��W ��EWLU�N/`8�`O�<ЁY��.7��p�Jo%^X���W���J�d�I��.�

�E��>Z�'wd�:%�]�]�6m�$�rb��[ځ�$����O���6E�SC�H���-k�BBv,���I��K��Œ�N �$ bb��>�a�#ʟ\�T%s��l�{�1~�ꎸBr��[t�i̤t$������ئ�_*u&��M�iOS��3-�[x��lp�+I񅌑bHO� ���/&Q���A��p"�HS2&ƫԶoFq���&"�t�niE�����u@��l(��Q�����`�a2�X�"w�/���=����ӡteK���3���k��N1|t�51� N�Cg|�~�]{�$�..��j�2&
�s��I��ȹ�`P�o���@��8�gQ�IOQeBTOX U��POus`���i��k₆=5�����b�L&��_	{(��,���-�Y5��4�y���D6%t��_I�/�Y�I�|7���]6� Xa<ѿ��J0A��EZ�����70F��a�1����>{���� ����[_�Ky�&�?>�O���ꩮ���6�g8�U�ۤ.�51c����0\�?��1�JΏ����OM��~�.�_�>	�+B8���Y{���N�66(�5��ͳR�C�F�ݾj�L�"�M\Y�`A�l����=.#��c�u2}	_Z�(��=� 	`��k�!�H&h�,�k�Ԣ�H"R%�SKfk�83qH���)A�u!���z#%��*��=CtTQ�]�Y�y`�y�=vvW�z�ʿ�V�Ŧ-I<�?�d������6�gm0k��`� d<"ج�LӃL��3���fэ�k����gG�ߤ*�H����I�.�C�em�;������_�q�}��6f���d����BŤ;%� Lo7�lq -�)�"5�Z�+	��&,���(iAM�/ห(���`s���Ҹ�F�<S[�v%cO���<p������H��E�����`(\�z= ����gI��9�K؂:�� �qR��J$`n��L[�n#��\���*L�]AH��2Lb��}o��g��]Ԡ������߻�P�f/��������26	��J���h��8gzՒ��?��J�;�,u;լ{�s<�9XDO��m]�킟:��*u�/�]�W��?� B,�e��qmԶu��W4�[�5��o�E�oRL#hL�:k���9�H��XBb���X����&HS&
>#1����f{�u�Y;J�2p5r=�0v������S�Ddg�a�G��ȗ���� zw���=��Ϫ8�j�0%Qmf�����"�w��������g8�b������"��+�(������`[0��a��-���֥���V���ѭ}=�f�F��3��#�v����\����ӎM��4c/��=k��9%?l�*�g�m�z(�Z]�B��g��!d3��9��\���}��h���=���s;�S��s���<Wt5DޖнWd�fw��e(3��kco�������o{H����q���h$���,��> �֣~�3_ǝg���S<uhf3�U+�1�
�qj�.0��z��/�&X�щ�n���l���Z�X��zi�ZL�x]���b>�i�)(J�@!����] ~�^I4���*j]���΄�~:�q/t��P4��dy�n��ɝX�ۅ�r���V���#au��,���Q��As��[_|0F��J?�k�9Ad%�:���N�CHq��]I��� �,�뢆$�д�(k_�+���� ��S_-8T�%8�N������5(Ak���u���,�� 3ZA��]|�D��X͉!��Bg�M�ۭ��.�sL d��i��3L�>�������rfzW#j���z	�p���!�KOFS��o�X����X����j��pF�[F/�mtYp�E�dm��B�<�E��+;Pq<F���$(�EP���ǒ�@��!9_)�{S+�~�В�3Jrm��tRy|�%����Q����	��#<�6���U꽑|9���Xs_KM�ô��2��V(&��k����_phceQL�p��8��Oqe�-�an� �3{_HsG!�N���y��8Pݫ�\�EzoF��2.S46e�@Tݭ�o�
#�ۀ���3�����y�ڰ4�q���K�u�QM]3C�r��?˪��'"��n��5��s�]9���{��r4��u\U�u3kw���9}[���ڒ�3��X�N.5;��l�)��13�J<��gD6R0��D���4|���S?A�KvC�����k���es-q�ޱ��ԭ���!�!�Suә��"t�O 潂?�4�/�F��!�'})�6�������e�P�1���7˩0����a���&.�P��۾S�}N/?��������̨"��b@b�=�V�~]P`������Ȝr�M���qaf�d���9 sǹ����/{�d�I��ּ^2�V�9��1N�R<�����5 3Fg����YnYq���x�Y�tS�������/_Յxk|%��=�W��$6W"6��4��tDS"��O�L^@C#^-�9�GT�8oj�#e�	���*�\�N8�XY&@�ݙ_ZY�NAهp�ܹ���n���h��˖�'��Vr�
�14h�fw�l�A�o����)u������3q<ͯ�\��d0jAxV/ߑ2�#��0��D����`ĉu�з�\���c�=_	�|=���n�~�6	Bw��]�N����sL~���.P���G��;��G���a0[�J4�j��2�(�ƶ���_��{�bA[+�+�_�����w��l�g��Jv��To�fۢ�
Xl��*�uJ	<�RW3�*�������
Z�Կ�/By�L��0����(�$�nfr��g��X����Ѫ��{Q|WJ�Kɣ�#DJ�B$H\�۩��m�UOY��!��p�3,�q���M�;��=�AT#7E��5ltrJm���Eo6ۯ�� ���' ���� �+��<��i R;��1�ZUE��%w9��H�5���$��Уv��nJ *��4�� ���_����>V���I2��Ā"TC�t��ǋ������!�;��T^օI{c�#��}�u]�-��v���砍�ET��j���$�1h�$�W�����L�L�Bt�y:�M�q��t�����Mx0Н�7�ٶ"�dO��K]E'�܏Ѫ�~�zoEs�? "ɦfӫH'���F��I�#�-~$��./mRI�1�+J,��HNq|⇧x����;|rW��o=f�++�j|5{�K��'mњBhڙ���ƈ�?��#H�6O%0��B��200�ɕ���w�eR���2I`�gsfPq+�!�cs����C9�,�hY�s�G��a���(|��J�-�����v�����u��ú\S�h#}$S�g��ҼN��|��V�V�j�c�h�O��"|{����p�x��H���5u�|������D鱎�����{gںSQ4���Vai�q�����F���A*V�^f����A�v�QL
+R>{3 2�XSB��4�e�t��I&kx5�p��\���y��A(Q������jI{�{r�d�o��f	�a�#���ֲ��@�r�N���!Ul��W�^�*��),�抰�����¾O�2�'k��������NS�����A4vo`�9Z�1{^�_&XU���H�M�	���\�)�l�PFP�7/N�4�n>
��]�,���w,��!,��͆�%뷛��IH��y눴܉��u����+=g����͡�>%��Š�-�SD���oq�uxVv+���(RM,u��Z>;}����ů���qg�m�Z9������_Mm�������i��5�k6�ߣ�X��ker�g�12[Q��5�bQqE�A��f�&���&u>� "������O���������mwD,��iP�ɧ.����Q��ڎ�
�a=U��=�T�s}�^0S�2���!�����-u��|�����I�$���fT�������;��tb�anCޘ#m��1�2 4.���_�ʋ��q.��ޞ����%����̺%ɔ-����.A���#�[�@�\�tΖ���)�OK�~�[�1��ei�s��Ţ�e�(��Iif{���֣�|�A�ۿr����@9� C¦N����4"�l�0�I���P�Ғv$�2���¥6x����rT� ���M���ל��S�h�Ի�����ɓu%����snz���4W�b�!��O�����LzUeE<�4O&QN)� b�� ��=�MK�a�% �Ǐ_�G[K�l�׮�/l!3r�s
Kɴ�&��x����B��9�i����=Q��2}�1���J�|����0�OMb���5�@ ��A���ppx[^@*��T�r��R�����3��]�����u\��YA� 6B�m��O��wv�>�~p�ÖB ��^��j7��,0��z̷(
����Hlt����Vg+�=��[�Ef*��x����~�5��ݞ2I>]p��/=�Q���*S���H�t3����{���#6ᢺ&hJ��˚� �mH4	��U�D��谦�$����&�eB�\�j;�2�a���}�D����d�R�'7�#J����dU4���,�j����9����o6�����?�e��JJҧ!eA[�w*���un9�F?oE�����Қ��}ߔ�tCr��Ў��ᩔ(������s���y���}��{�Uw�;����'���~�*�h�v���b�) ��\���q�S����՝N:!�fu�\����cY�H�E��G��_��{hx���"=N�s��v�bƱu*O�w�Ƥ֧�x�	�F���@������nX^�E�U�x�6����Ĝ�NYw���@�r�[�X]gpϤ�����~}atV�A@�\]^ ��7��/�%��F`���u�I�9)���,�	�:e*��O2ͦ3��7�	础A�16��i	O�3&��'/O�Xc�W���L��:�gM9��	���Q��L&9?-�x�'�;�Ţ}�dT4�,��>W��x�h�j������fs����n.�b2�<�$'�r�a̒�x� Я;Ty:�	9p��0(�5���r�9�-V�C�i��I���������_�E���ѥ�Mؾ��D��,qڅ<V������;q�L�����Y�98Cӎ�Je�'��õ�.�[V�DG^/[��L��lT3�O�n|��'��Wk����~�m
�ڇ�w���-c��-�=��a��g�?�А�F�N��a��.�T�l��3a�$�{��c�4K��=���^F-rcVl#�IN�d��/f�߃�#�k��I���l@����\�l�5�[�[L̻��R)�����/;upܙ�C���mk�Y���$����x�E�)�',������R��)�X�fM��qdw&��}0��e9+��y��|G��ujq�f�8f��5Nl��|E�$��%�E�sS[\ʵ�C/�֩�/ĹT�[����k-*�詺��	*�y�7*s�K����[��_!����Ox2��4u��_I�o� KMT��,]�fď�?����6���2^�� ^]���`��r!T�I�l��/��˖Wz��J%e��-!-릤)��˼R����6\�Z�'���"��������D�s��zeM�?��FWW����*��3P*	�,d�-}�6�( 1u<>�mɭ}Z�^��A�-��4D�J�B�6 ��N��Z�{#�pך��}f�[K�!�	�����irh�(�oT��{����&����2.�p|U�R���0�n2�{�9�I�o��T0���CQ<��������Y$�"�&`�sA{*5DBܲ��֩XB�?�"���{�waU��౏XC�G���K��c�0Pe����.�	�'aC(�)�/�N�a')���I�y	_v0�[���EWv�c��weQxF+U��H,	*<�,x'�*��*�1�?�l��q�;O^��P�׿��PE���p�p�vw8�`酨�-��^7n*��!��!����/��$�5F��0It���9���Cl/��i7�
g�2�zN=�oa,9�`V���G�T(�J�҂7{[�B�W#�E�I�>ٛ��:�癥3�Rc��*H�!W��AlnbL>�c�_4��sCQ�V���w�p� #�T�&����	�������'������ޔ�� J٢�A���{"2d��M�tSe�R���ɇ+qn�iD�y�*��'#�����[�_:u�PS���U�"��y+�B~W	��BL�U�o����������_(�a!�QULI���B�|������2 �;|��}��z͐7] T�Q`�#�Z����Qi��<������y���(���ѩp�ռˈO�&�w��݆ $���<�pQ���k/YS
n��T�����l�%Ca�C�g�;�6(i�`��ZY���\c����M�`S�W�g͹`�ʺZ�O�@�B�:ڝhN��8$�H���Cf(�Z0��<"�3^*��-����/f�.�/U:��iT(��z��e{6�w�!�)�U�&1��B��,P���ˏ���弖1�*yps����{͕aFV�B�$�t���c��Z`?�KΝdv �)�����L��壧�Y桞���x��n�%#sC�t�����Z>�濶Y(���S�^/��.=QC[��
��~=���^�պ{_�H;i�^��i8�c���Y��C:��]+b���g�}_���#�H��聰ص�:5�����V�Uk�CU�;��p+�@�"���pحb2L�	�|7�27�V�Y����
k�ےR�L��o����n:� H5��ԃ�0�V��o�}ַ��R�h��.��0\v��\�`��?8�y�N���R��٬�)K���h+$ y�4�y��/�פ��X�kx;B)A�Ζ�E��y)A�����IqF[�$-�O��3>����0�%�<��V��c"|�񰱪)���
�]z� /ޯMAڽ���Y(I|��F7�Vg��0 
�U#�P2\A���e�	<R��heJq��JB�0�@�MW[1>��!��9���Je�'|<j����3yx8���%�\�i �q��m�"��>P�"�v"�-V��?��wc����J3���J�J�eh<-c����T��=բ37��G��si"s��^���*���UN~=��IF�࿪��K��wg,���p��f �Y!�bpk�4�2��$7p���"�T����� *u�؃<sF�g}��!p7"N2r�S}�U[�L+1�Sm�����2�����-&��d��w>�mx�6�����E�nOT�=���z?����������R�8�_����-zsN2e=⤒I�j��8Xx=��l#I����l�lN\�vQ��	�p�������������^#_��[����SBf�I^�:����%�Vu�(��.��8���hrs���# ��&���+�E�
�mw~�tG�4ɅM�;;fm6*��oɎe��Z�Y�A9���5�_�����5�áR�p�T ���T�y�������6��)M�rZRm�44�ٛ�l��E����ǩ]�M˺C� �끩KK5��U�a6v3�tC�״��>����`�I��]nE�)�ƉV�j�/�gR4�,��n��񴽿�ț{J"TƓ?y�������(���Uۑ�jOc*��T��j�LT@$_X��Ea���n&�}_��LԞ�6�]�����}��g���ϟ�^�AdrcQs��k9Z��d
�w�F��u�Uj닷����wT/�LtQ��_"�B,���	-�#��>�#�X�Bf��*,��Ɵ8�E\�UD��蝜^Ǆ�*�����(��!�4<�m��u��&E��?C� ��XZ4��b�8B�k����� ��;;o�!q���*�$�����NW{t@�M�Z�'�.d��g��j������nK�1"EV@t��I�㰱}�,ܶHR`X�т�@H3:���NE�4=��5WJ�s=��p��?��,=�6)0��ꦆ<=�5�D���m<�1
��yO�YH���N#}��ƒ� ��|���ԚWp�/����v/���!}�;����|� r��M��/�t��I/���98�����ڡ�w��r��J�8��`���#�Av<�Y�9+���%QW�c�h�#v� �ɋ��u�,/[�P[���;?/`*b��M���2�\����eU��2$��@	�\{ӕ�:��Ho�&��g$��{r5�q�Xh��)��F�?�1���D�uc�b����ap)�l���vd�L���PN1�h����b*O��>�٪﷫ߣ�Ҩ���J�B�f�~���T9GM���=e��w�r@�'�DF�A3�[����6��R����:���˓6�f� /��k ����3��g��}��Y!��*7����Z�G"����� �}�f�A�h�4j꨾]bݝ���uRd_z$�2��A{ߧ��>M�_Z���\?3оg]$.�
I������J4$�_�we�͛�"�;��[���e�
`NW����Ʌo��p��E3��:���SF|Q�g�J6�<d�ϱ�����6h�z�C�O�K�p�ؑ\;I��:�?�bxw�h���;4�p��m�2�3�F��}�]ֹ�E�Pq������O�6�DB:$?�X��ӯ��;�x)G��)\i6u48C��"e��<n����>��!
H6��_��}�_#��|% ���6�a~|S���;R{��4��Y�K�􎱢����e���s�;e�`���p?DJp)P����y�3�l���J�����#��tb1F�.�E�j��yۣP�c���Y��{o� �aI�����la5d���-]A
_��]�lL��6}��~��z�ф|-z���^��v�9��4�i]#����NRJ�,��hh���LI5�mܾ6@>���j�����K�t��X�z2i�l��j��t���b�u �p�ZF���"h���X%G��d�{�f���e2ka��wǡ�l���!��*�u���8-�p�0E�5������W^�&���A���&��1�]����>v;�o�<���_X�5@��n��<ei���ѻU��m���7�<W;ѯ͡3=�B���@�yr���>��.��+[E
�?ٟ�y?Q������邺&�����|-F<�%�T��pi�ˠX��+|��_�G�^��Z h�LS�-�)Mml'*]�[��Y���\O�4Sq�Vo��d2��(TS��(v �}o��i��gbx�@�z��o=�F�'�;�E�Tl����Ϗr�QeH���o���>Мu��\�)�C�H�
���`\�a{�E��~k���\##]� L&��,4.�~�Ő>E�u5;���+���G_�ҙ�� �w��M����S?�E>� "u��ǟ]7��:�d��"x�yQq�7�p�3J���ə��u���ج��qω���3X�|9�E�B��{��d��"�i�JY��G�M$K� -f��j�[Xg#��F�� �	Wj���t�H�0�ri�q���|C�[��>-�Cw��H2/����M淠�+�ǳ�flzO�.`Ã>�P	�:υ�P���|ć�O�rV��4.(�Iȴ��%9N����� p�M�yr��\~\�驐�P�V*
�m�'�vw�l�?X���!+)�.. �uc��'�s�Y@陟H�=�u\��JJ���E�(�
�"�yL,�P�}s�G9�X
5���{�z�U��3UJ���%�8W��ǅ�V]�X~إh 
���a(�_;)2�Ӊ�-��~�dqa\�1<�z���Ygc��g=y\������u�=�D��[�P{�A��I�|{݈横ejhĶV^Q���9���qed�ԉu��qz�ḉ���ɾ}��� �jP�<�!P=�m�³�L"�r��%�?�Z��y�z�1�(�Px��e��P�,
��F[�!?2�:s��ǟ�����������iKU��!d�n��X&��
w�����F��DX��{Ԁbgo�u�SK6��M<�<�����X"a#iӵ$�W�6RxK�F��8[�B┇�A�[{��|L0h'�N?��ѣ��%�~Z��G�c�i��n~5J��Qp41Q�ܛ�����l��^ѤU����{}�2�%г�҄�P���4�Y�X@�U{&'
 �KK���@4���L�>WJv}�e�v�znV��YM��r�窹1�Q�� &O�j9>���h�!�@���)/Bx *��@��4�=�è~P�\��Ĥs�3�͵)t���<&��� D�Xb�"���U뼦��V���$��OD ��-�����/rjD��$i�+��}v�ȭ�#�7�8G�H��~[�G�����I��dE:��ڼ(Q�����Ք~3+ p�"T����
�d�� z�2���jW�ݨ��x��4{`��Y�KE�I�FC7������˝��5�Tw��V�XJ��O8�&�d�9�f��b���r�|w,���#�a��J�ڼe�nC�zq��Aq���UݑBJ���n�(�x�d��K�3��W������	\��ٗ������r&s����G����g%xW�O�`�a�-pP�g]�dWA�ռs�q��n+^!1`2g)�����5U�hb�:ɚ�/��*�ݐ��d�Se�Qt�_�?ث���Hۭ`�d���ʽ� 4-��T�Ok������k����V�d=�p�G0�&`���=�t�a��Ͽ�eV�Tʮ5����BI\聨�WBy$r��c��o��/T5�ow~�Q��t]@(�A��|m:Ȟ�α���ioLѳ�	϶��>L���c��sk0�����@���u��/�h᝜���U�YH�/Z(V�+�8n
訯�@r�{q�<�����TAy�F�;ᐖ	��l�3��y�����k��0��4�E���{�w������1�x�\Om��xΠ���i��A+aC/Ov�!�+?��AM@~bó�E�_���EVn��������� ��I��A��NJl���OY]� �)R��68�X�U����v.��� �X���P�n�7���N��%��[V_)������0��БX�uM�Q��H�vh�'U��z��8(T�z�*���FӮ������l��.��
>Rsx�V�E[gV��ȟ�y�>���5ׇ�gTr:�J���Lh����{H�R�4ÙX��,lB�i�w	V��LS�ע�E������ݼ�>���԰���Bn*�C7K.;�`����QLq���
T� �Cl�l}��:G|��.��(	a�3���4�h��P��!m��iD�^�Ë�i�����0ӝ/��p; ?3ѭ�8��qģ�5�'/��es��N=��.�1�j�e7��պ̦�����"�O�m��՟���<K�� �Lc��{�V�E׀9W�2��"`�#��uy�\Ew`eE�e8��X	d����)zDM8�L�� Y�~��6��u+@!�J �j��&���p�l�lK��$�X��cS�Rr�;����|��(�.�
a�m��YX��Si��H#L�p.��#T�I\�F�I�s�w�^�ԯZ~B6�As��kŝe����C7#��:��k�w�(UC��*��>m�dP.�+:�РL99����ܖ�X��j���U�g7�[�{)�i���|�cG�4�u��>�>�`�F��,zo�!�;�d^|#�{'�H�.������!R�9"����Ok�j4�8���wA���������J�V]^�NJ��=8�\�� /�5q.�Adο�{�J~���`:ߔ��,*2���/'������tl��A6����T��p.�Ə�R*��Xb$��49Hkdu���Fcu���X_���dfc���.62��5�R���0��y����z_6�R{�v�+RZQ����-��C��ت�\���Fieu�6z� o�0��~�1'�y��T��&$�����œ�c7YWӈ���A�����7��uR�2�Ɇ�-�,��~$hp_�� ��Z 4���;^�l���+.��E%�/�V!쿩-�[�P�"aQ-��̨�O�*��c%��a?��C~'�
v����b_�:C�����y�M�����oi�hg�<)����e�6(���X����cQ���hN����$����e��^F�3<��*QH
�_�����KBU��e�ۖ��3�3���Do78¨C��',d��	鶐���V�nW�O��ZS�
���e�d��[�@6�J� ��Tԗ�W���Y/^��Y��&S��JukUGB޵(�*h�G��7�)��:��"��uy1��1	#��Lׅ滼,���+�|TZH���|��#lʥ����U�|���4+׎l�sfј�%�m�z�i��l@��(9���#�^��h{W18�o*�8�x�o8ߔS�����i(xV�S�AVBrz�u&ʺ�����2�o���t)�����U�+�E���3�#�n�WX��LkG}�L�D�`�Pr��r�bvzU���*�Z�o�0�є��;�Kz=r���i�y�m�3o@�@;t��W>|l��s��޲z���Up���Hj��Um6���I4Ǡ�9�Xַ���d4t��;�k�� 
�� �D�ɒ`�ܜ�}��R�&�j����R��'�2����`�e�mXP�s���p�P�/[��x.�Lp�=�u�悷a�֜�`�qr��#Љ�����0����}ǎ�5�|����E1q_uj�E0wJ��xAs���j��[Çܳ���0Ǖ�9�6�5�PP�V���b\[����ڼu��IW_��Hu�B�6�m*���Q��7��ͬ����]V��z�'�,-o0�\���(%Gr��<غ��3����!�ٕX�(L�K}���1���Y��*�'t������37�&_�Tc}�N�F%��=IŅ{T�Ԛ�vN����u�}�L��B[5��뉔7,��{7�ך�DO�s���H�ۇ��
����q~�;�ׇ��iC�E�}+�t\H������]*"X�oZ&����9zw���ڟn�uV7����#EC1Ϣ\���dy�:�ޙr&����ض�`t"��6��9x8>�@����1����p�a�?,ܙB�k��;4&��(�8�-����-���{D�щaBH�����Y����}��� O�h�p�ߖ�����ڰg�w��oc'��hӻ�R��C�Yw�5�p�u+��/�Ĉm�6}5��J�`4�Rl���U1	}��������>
��}�7���J\M��MַR����b�1bc��:k��i��s5�!b��_�w��G�r��^%"S}��9��V�O� �[R^lus�Ql[�V6<���T[��γT����CNUL�CX����?|��ĊU�v��9h*��`�	���}�eC͵� �Ԏ6�v��
U4��z�6��x�=U�ʶ�Ө���M�!�ů�oBy�.��vK)�7�����^�S%
������j)6�{���^�����m	�p`���d�تK�2��(y�)x���V�q�Z}!����$�S���i17��Y�\ ��4�F�6	����{fj�t���M���W��+��z5&(җ��z�>�Lg����蔐[���&q6���o<۵*P^eF�=���}���m�+���\"$���D�
�1iRz�)>�fk�4����tŕ�z<��	��߻��)?��hLw^�G�O�h� 3%���<��4��I�2s����
��EcӐM�;��QE��qC�ۨp�H���
�?o�"�@ �PiV �"ǁ��;L���u"<OG����˂(O�k�2��9�譗V�"���dp��$�f
?����KPB@���/A�bș9�D��z[�	 S�_Mbv�w�"	2x���|F�n���2�~���T����W�-d�f�~9�l��Ȉ�^�c�]��_�q���-�'kJ?Dk�W-)b�$u[X���l�\��� y�yV0\��:�)�K����qž�[���i��L�5�"�q�a���g$�fU�!��� 8��N�RGTJ?=��sL�r�V:�Sg��T�����,��Z�C�2эKz[�m5��|�sC͔<n"�"�6:�P3j̠H8z�N�ti�q��>f�y���ㆰ�}�Xc�k�S�����?�~a�t<}S���� :������J΋>~��R�窱k�
��R�{�}L����Ny�J�\�+K2�w�kГ��ʷ�S��4P:"�:P��JJ������k0�͔U��T��ՀÀ�6}X���ȓI��,�#�ϸ����K���ˇ��2�/���y4J�%&�˪Z�ԩE�8�Op�G=��X�A�kd*��I�o�uѓ�rt.u�z6g12�҄�D0�?���
;"��ҡ�9.J�U�3'��		W=$'�T��<��KT�69E	��Z�Kta�ϋ�{�pq�{�~�hIl����bdK���@�2^�����4�g��s50܄G+�<�O�����Z�YN���O�]�����X9�'(�;@Fr����r��}3��Y�?���n|�>�R�g_Ly�����~\�)�.�H�'Y����g���x&,X�~���ޢ�/����E1��d�F��gRȈ�N���*�6k�B���;2/p�*7����	�#5�&�����Q��L6/�+p�F�/�s#*��S�K��w�,��+�.� r�r͟�:���X���㥃�
�{���T|h����'�X��V�;�MX��
vd2_�挍��,�p�P�;}�t�=��0�}�-�T�óg$-��f�װ#Ss����B�6����Ҳ�5�C��bCf�L���Ç�c��"�X�.څ�{<�jd3�b���q=EF�;���I'ͮ?�4פ�8�/,�	��F��E͙��CȏӖ��X$=���ǊF�W�3���q�ؠ^ �K�.���(��Ba�Nsx'q�C%��2�s��:�^"*��H��p�W34Xf,�:m4����	����F �Υ\�[��9Cj��AU�}d�+�Z��4Z�2�aӚI6��=ÚZ9�d�^b����״��!n==�, ����7z�z�҈�ML�n���Z1־n!��:��=�A)�C���3`��7fO��#���˓$��ٰ@�"}vݖg(�����jc�@�U��=��"CJ)��o�	4fD�I���|8� ���=-;�x�l<2���F����O�����%� ��&A��f������d�����=j�X�����)���������.�)w~���f0W�����k�_�^HLG��/�]1?�6�@��1FIik��nz&�K.r�'�7J�mD,�`g������$�ٸ��4�dx�9i�4o�gNm�%ٶ��F͙����G �0*���Թ�,5
�/oj����G��/��EV�8�O�@۲.#�;�R����Þ���\�ݣ�>C�U�ݎ��$�[FE9��`l�\�@x��1�!�#��X�mh���R�*"�t���'�)P��c��#ܠ)�o�zW*��q�a� &Wa�,̂^ � ����?�+��4�8'zbN�Y�z�>w���ƙ ��MT�	~�H����=��˖#��_��<kÓC"��y��eF@���F��"AR��u#=i����;�G�h�O����_���թ�� �8�#��D>5������;3&�CT�F8r�.���n��B�"���\���T����a3�M��9�s�f_7%���ᡦ)��N�i��a�1�E��`�n=Fx7�������h�Y7�i#�5+�� mJ����!�v	q�? CÈ��ܓ"�l�f(3�����E���M\��cK��
�~�	��/�_[h{D�T+���a�,�`��Н<�e5��U�����_���6�+�,���Jr�V�n�* ��wz�aD����mX:������*G+�V6c7�U/�w��@�;I�Ҳ �y���N���d�+u��Ӗb��,�CB���Z@�	�7�`C��X�}�����3;	�Ƹ��ƽ�x�	��Q]9����pCH#�؀r���]c�A�o�ކ~UM*���U�p��f��a-�n�,8��tn��L��GF�C,M,���~n��S4�2�+�k��]�A����9�e�p_:S��)u�A����#(�<�a%���tΫ�K�z�X�g_B�Uyg���П���k>�[�DSo�`�9�0����3J�$=�+�x��f�Դ48Ҩ[򴾾죗���*���>x��Q稙/��ܤ��2JK�v.��w���%\�[���'r�0k��=荂�\�>4�YEL���(ozeX�w`ٛ�ٻv� 9�'h�ؐ(�h��s�ǭ!�[��4qc��꽳!���c:?�-kA]�̼D!�a�2Vu�F��nm���@����KV�e
y�5��?�CqC�� �,I)�$�}؃��"�iFǔ�5�,���>2� 0g��s8�"��)'�
�=!K^D�!@ٹiQ�`p"T}l�J��Qmd�z�dW�wb�'�s7�����}� �Յ��,"<W�������y�D�=>����>��@9�S�������#����>���cQRჀ�m�LЍ���	��;�}�	b��e��F�Zg�{���{]�7��z��|�@��|߻Q��6'^���k��_M����iU�=F����'��>f�<0�Sp�[D<u�MeJ�q�=;S���o���iԙ��wh^^�O���2���uD|%���L��C�O�	 �L���5L��Ĵ��a��Vg�u�����I �ul$��_�����(��k�֔�s"b�bvh=�|����)�#�"y���}1̍�O���^X8���x��	�_��a�z���|;z����`<��4�%��O �j���UF�o�a�����d��L�3韕�T��>�����Ouf���-�*�8���5 Dz��Ge�e<�J��9�FX�-�}HlRdb���)��z����R��f/�u#+�P��Za�e���z�DG7�Z]�x�w�l��hU��43iEXрBCVN�nA��Ŝ�61�WG�!�_%[P�b�Mf51��h�o��X����H����
�
V�8�+��/�1�F�7Uc���]�q�����-�U��꧞߽�*���<}����[�n��mq���J�����M/:�l�w.Y���"�a燅}Q�	k�����o����8�1M�׍;p�8wE
�ڹ�R9��C�IGY_��a�M���0���>�S�L�"�ig���D��j�\��rԵ�0�J��Bv��[�b��KbI���!��Ze���|c����F�h7N�^qg��k.�Q��A�a��39-V�(�e�\Ï�bR*��U���BJ*4Ї�� �ã&��˽0�X�Β3�ɐa{Bs��V�n�H��:�:J�K��\}C�}�`���e��L;y��|N�R!K�h�t	��xЂ�)����&�n�7iK?]U(��ø��꼘i4��ЏȻ���b�����&E`Z���c!�A}pJ��a��Mu����k;N�CA�=e�.j��ک\�*]�\���,N�Zm�Q��t�#���,ZG��A�V�T��/J</�mp&˶M�����g"3.�xc垮�h����[�텏��"1JQ��w�j�Qӫ;�[782h�v�� UT����a\9�4{EІEQ`���|��U�Sݍ���X��=�yn;=va�6A�ܕG��Y�����$b�pc?1p��tj���QuM��+U^+\�f����Gm�B�w�&����Cz�ly��E����H�)E�x�H����o���i�P4��D>n��`��Ü�ゃ�\i2ɱ�Up���F��:��r]s�4F�O#��B��RD��='��r/��+#�k@�L��� Z�}�M�&��3�5�׫��B5R�j&A�%{?_�O����Q�;�_N(���OK�� %k�w6��iv���>�� ���-��9A� `c��@Q+Ǭ�����"��N�9U��,��vN���L��- �ҋ�_.x�;��u^���!��$�Nӓ�>���ļG�.��5�f:Nf���Yh�a= �Y�� Fa�	��ɯ�."���= �V<�9�� `>��T�c�L��7�F'Y`�O��j�f��|��Ϛ���"���y��:���?(9���4�H﹚�',/�J���7��97��|�'�ś[ ���B����7�R��S2�9rdR։���羼��U%(w�CG_���^���Z-��ָ�Q	FJ\w��Du�gu�,�5�T6��?� �k��KI�*��<�$>kc�� �]��w��KX��|!�~�'��5=��-�w��i���K��7�(1�_�W?�;)$?��!��a
�J��=�T*��Y��a3��M�}]��Imd�w�����ͺ���WH��M[��X�|�Rs��g�*I��
}��<�3�X�c�ÿ�`�'����H�����b1�j�u���`5�u���ݕpf��+�Nw=���|�6���Q2=p�3��<�v��b���5������V�GF��%�UD�|c/X]+����0D��p��t �N����܀9�r������'5����\s<��+���y~��sl1�ܱ~g�`�@�^�0��F�;���ݤXK]o�3���D �����
%������Q��3o���������l�/���&j	�
�3Y�� ��ppt"�-�9k�E?�Ndz.fC��0���D�zG�EfX�|��%�%]S.� D�I�W���_����F;����:X�Uۍ[�A��:j�|A���_�D�g	�&���m?I/.R��b�C��dW�e*���u�h�,���੺����N<�ko�����tO�M��v;D���q��"I$�e�=�@�my	���G���1��M�6��K`��$�L^�-c�h�<�2����N�~g|1n���-<���(ڴ_��e���
 �D_ӝ"������ko�_e C{��8yO��.��� 7�~���o��~&:��މ���c���|�B��>����@ī%N���
-*�x�:�k�m�<ݻ�ED�����1���1G�1q�V���U_���1]�nu,GJ����ʰk�d�n������z2��X�rSɕ.ݥ�N����QZa.�[씧Z�#L�z�f�ui.`��M�6���z��|�x2���V^�8 �W�Nu�i`蘱�ѫm;�DY����U���h��)����"]F=]F_� ��V���1��|ɯ����8�<E&�!�
��;6=�Y����Tq�����I�8�`���O��LM�$W�թk��]5 �w��-o6�q~.��}�i�2��?����[��
��[�_�6i��]�{� &�o�
�ơN����v�ݰ�������}0?�m�U���7����s<o��X�����]\�~�6o�9ze�x���,ׯ�sY��?.�"T�����|TL���^� �e����8�Ec�悽�O)̮1K�y?0�]�Ɍ{P��u�}LI���Tw�1<u^nl�4�WA�y��[�}{V�`�y{n,�"foQ��𤐨�>�g0@�V�*���Y��Q	f�����_͢<��8������?�F�h#��G4K�n�q�F�=!���h�[H�����"��y�?�K�qi\c�s�J�@ԙ8�6&�"�MC��̯`dɘTa�ϛ�C������֘.�����M�� G��+P=5�9�2���7�m��i(�>l�);<���ʯ(J����*��iD|N,�ͻ�2d�8]�(Qv���.n7�2��H��%���i����@���=�鏻�9�6=��ru��;��6�6�SM�n���o�)_t�Ȃ��{��Ш�B!��j�h���e�0)SXR+TŘ4�p�0p�� A�f��3��z	91	.��{?@CM�U���py�[1�wL�7���$5����\I���!C��Lr��|�6�wq�|hQ�}�M�rʉ6��v)X	��#��S������s���̐����/S���ջ�1#AS�o�o�}��GT��&�dr֞b�֨9<A���b:u �+~c�a�����pr(ֻ"��v�R�Ȩ*�OVo�1����Z��ʠ0�_��pXSM���}�K/U��	R���ϐD�8��u������bC��%�OT��}���cw%JT	�ǃ�
d ��ȸ2�jv.+fki0(̸H���¼�����"��" �9�O�&���l��.^�Y_xq|�%�PVX8����n��,B�z�B�Kb���X�;A}�C�)F/�.�Y��C4����.�	%}̿�r�H�9��&��{ݧ����nb*�9l��5��Q#l�+���D�~��b��5Z���ZgW���Ў��� A]�����z:����,�2(c2ub4�!�M�����,��8�""M�HIPM�t�/i'^ɥ؃�n�+�#��smL��E?�!�N���M���)C�ZFКh�kw ]F:ϸ��z�x�fL�1��J��D�3����5T_Q	!�:M鷌ے�j���EB=}�l�T���=���^v�H���mJ���_z0��;n�js�l;��!�r��0+�h�����?�x������B�t��9o$~;���kV��7�,ԴY�.	� ���v����y�i�k��!Y17�vFe��[�<�{��P�I��궖:|�:�
��b����5��=)`�&�M���ɤ���W��$YK� ?�&��)7�1;�J��^y���/]rʚ�@�]�h��e��l!����fe��m���\K .C8:i�)rb�������.��`�8(ʙ�� �<`fa��|7E	ϛ}j]b�S�^����zK��P45���t�Ŕ�xF9>lr{��&�MX����LC��S����)��v˅�
b.�s$�ƾV;Þ��-
���S�v�a�ƶM���e(oXIha�0ߐi��$�FI�ف�_捹��[�]֐p2� Z+�v��RJ��͖�����q� !LƍE�[���ީ�Q@�Nі[��}� '��>�^<��*�PqQ�]{ëm�04'H���Xa���v�p���:�gvӜ�N�v�j�n?���reL1�_{.�C	��.�؉���F����w�$�*�T�a�{�b��N��#��^f����"��P��f�!��7@hx�w�Ӕh��v�[2j�N�~I-�ς"�����G;2�^���oE��Q+�e�tP��֢cL�3����<v����y���γhDW�7r2���1^3,�	#/�sH�]>C���K!��B2~ɪ h�Ĵ�5R���ȯ7��W/�&�þ�q?JA�n}���{�7�C�A���-�k�k�	I�Ǘa�<b���'h�$)���t�F��öhd}�(>��}QT,�b�){�.�h�� W
D4ѐ:�$�`.���5�r��á:Ɵ�C^���Ѵ5�m�O`]�h1H:<���^�]zAЊ�M4=(�j�IɥA�jb8n�"9m�5�)�p�@_�c��5�˵���w�2�*��/��,��;�j�bJL�j���aגE��<z�!��*�� �O��]�;#|è3� Ŏ���r��N�p��7c�����8i�'���O�T�>�\�b!�pc��A��k���
X�Д0��Od���j�5Zn	}xm����*�����1����� W	�8����y��S�v�+,�{�1��ص��~�R��hN��ev���]ys��*�J�Z�X�E@W�vO1�ɄT)22�N��P{ճ[�Y$��D#h8��9VW>����Z(�]积H�}���4�(PlN�����d"+�����p��-r��
A2>[���J��Ͽ�ɚ'g�e�Fg~v�y��e��&�)Hᕫ�q�g�^��s�U�&[�0v�>(%Ѿ$a�sS�l�2q�}q���4(�>� �4E��v�m'��4�p�:$�x��r�l��[x���_��9J���
�*V e������$���^���!%g<ST(w��t�EY��дx^�`��}m��Ę�ӄN�m��ۯ�9�O�a��r�����j���X�!>7^u�x�y�䥇eN�e�!85435Z�}>A����:/��u�3����5�ᝌR�H�H`	�,ԬG޶H?s�����T�}/�f/��Rt;��@P�������������&�jä��kH��'ߘ6���jH�.�-LΚ�ح�u�W���5�x?�BHi���i��	�Jp�[��v���g�n��D�L�`f�n�4�� W(AP�n��[�wZ��$�\�������b����T�G����d�����}�E�(`f;`���z&*����잿8�Lk�KT�l��K�.�fek�)ts����Bgʴ�6��	X[t�xG�m.��S��f-n�j��yH�I!^��t����H����*-���\-v�dPu�J��<ua-~���p�������|{%����S�%O}�:>E��h�v ��9>;4�ih���)���8��~����	�",�g��C��U��w�Z��)�'0[��09�Ez�o�o��H}�������fɍ�2v
�̭��e�v}	�[������&�,�t�'?�#�p)���r�b�v�S��.��ZqCi"Eo���-�8���$��t$�*Z��Zo6�4�cV��E,Ys��C��@�\7�/pI��h���#ʃ�&mT���Uf���lJ���G�U�-`��г�!R�Ĵ~`�0�Ce"�tc���<���%��c<���U%.\�v���ڏϟ��Y�
��S%g�r�Ai�uT�B*Q霛*E���k0��M�����?U�v+��f�`5�Z*�k�zHh��I�BPPG5��<�GȖ�'�7�̷@+.��9ڋ�:�]����t0�/]�~��*�@�[��#�2��7,WT��Rcqz�M�uDar&	��>�$�����sj-�8����2��>�;�]�G(ǫӿ�a���P�j�Vr�<�Q�3>,a���xsr���Pe�V�F$���B�m�+q���:�Y�<����sV����Dhl��~��/��G�Б��y�{�;�b���Z���H�1(�j&����!,�D+YT3װ�ݤk׀w����+)�J�>鵑���x�������l�R��Es�v+�;�J�~��QW�K�*5�L.����oU��n�|�����׊%�}���	ZU-��5�4 �w���WDrp}AA2"�����<��$����+�a�Lu~Y1Y�ak�����O���{O�/��*�M�L���J�1{��N�.#���Y�P9�^OdVb|~�Pw����ۓ��B�C�sy;�v`"o�sYic��7r�w�0���0̛Ƣߑ�kv���I�|�h�D�8��}��Hmz�e�7�m�7D�m���h��V_�&�p�BU)z�H�hD���#DE�G�����tK�e`���]��o�.Hg���p�׮�{$�W���  �����18·*�ϊ�Da�������N�[�D[&�5����ҽ//p�q�j�A����3�b�[/���mp�ThÈI��os�����0�~�d��p�����5��]�YPa�m;B����"L{��	Ê����?߂���C|�B��qIV7�V�/��.�ҷ�F��S���|c��,�>գ�T=�&�5=2����-S� �9���k �d����+v�#~u�G��3���f'@f�T�l��F��� �m���8�.�)��*��@$IB��hZ��,�w2jk�/���\��� ?��C-���0L�} �[���9Bn�F��&���8�Q� c-������j�I�wO{��N\��h��F�:��}�C���x�u�1���'21ɤ&J��U��ݍb��m�N�=�G:T4����R�����kyB��f�n��� �[�|u��e�n��ʻ� JNt�i��wT�*y!CE2sY�;�ZWWf�v�P8S�
�(2����m��Z^
�Eѿ����:a���F\3��]`�(g&*�}�E�lTc��ݫ^Nl 
�i�9��;zX+�=�އuH����Hxl��&_����]��'�����niz%��1��x��%$��'����M�#f7��WH��EG�/[#���)�֢��ZZUO�ASx���6��y�b�-��r��g�l��s��T�$��/���0Y�D'pX�*����3 �׭r�z�|c�noZF���7�gSS�rD� $�[��G�A�A��h�B��ޜ�ި�l��J&ud��6ipW���d �*�Rn�-2K�����d&���N5����A��1"9�P�������G�Flp�[h+�~R<�ڮ�T���?Εu��?װ�5Ksy TwY�?@����h�2+W�,�@ѸYi�Y��$F=��0:"H0E��$�zʖ�)!�ϊ����Cg�9���+����]���b�~P��9�U`�U�h�?2��g"����cֵ��>��Ԅ):�d\N)f��u�U"�8!�1��'����X��j����|$�
N���b�"'�neF�f"�����7n9_*�7+ܯ���7��R�t�� i��d�^��p�ˏH�e�^��C���XH�h����`$p��&�lI�!n�e59�0���|s����ɊȦ��'���j�F�զ����ӬIF��;��,�ش/�v���yu�r�h��P���8�'%qB��@:cu��D����Ў
�G"�m8��m2�91���Ĳk���%*��NP��V:a�q=tb��m�j����G����Q�Z[Z;�=�Gx�4Q8�������8�k�8�[lo�!�"��Z����x8�Qǈ��I�q�)x��#EXK+_�;M���2Z�~�Q$���]��쉆�K�I�TJ��G�訋��s�qQ�Idm�C���/_�`Ԕe��?��c��re�<D_����SJ߻�}�1g��ޢ�������uLLϲ�Y,�mܐ��2m��{(���O7�6x�f�z����N�9� j2�H�@���<��Soq�$��I�+!�X�+�j[�ɽ(�U�eY�C1�oly:��8p�ڍc�=��<�=��ĝ5����6��N�f)2�x,�𳩰�(�Lh�ƅ2��p
u&Mv�̍w���)�]�*��fr�c��f܋̾��C��	5�?0���y��d�;	��T�ޙNK[{r$�'�~W6PO��p�����!w�:��M��'��-2��[�rR�J�B�N4H� ��譏6+ ��FG��	H�	[�V�=l��?0��	�%����%B�Bh���>K?$F�+��dQ6�-�����~`��ϩ~�_ۄG�y��A�� UK:�c(5�ڷ�^��L3�y�K=Or�L�'Fߪ��z��E���m�`�N���&G�F)5�=��I�'ݨ�ȝ�^����� J$���rnQh/r	GԶ�$�/�l#�5-��ɑ/_��
a�Ob������9y�D�*�\,�s�H!XOxV��y3��<ƺ�s�u�����3�	�
�ݗ��/��Q��'�S��J�7�L�N=hn��̶I#f�|��U�^.�Y�_�]͛z�K��5��=ro�Y
�Ny�q��D/K��ED��"�@�%��Q�"?�N3F4���>ئ�;�ViI�|�p���y%Ƴ���f9��������D|BTC{�`E29"�K��Q��ɸoR%����ը<�es�<r1?�W+$y�'�,���K�8ü;��ȜӦ��U)V�(@l�[z8門y >5��^��TCb���d-=���L�T?�	�����_�D��q�YσƦ�y�5��V2�6���CL�J��`uř��������W+/1-O�u��~	��Z,�4�@��O�b�AU=�c~Pk�^ӂJWE\7e5]t�:��X�����d!��.�0�p�(� 9����+�����p'.�\	[l)mA<J~V"(�֛٬�[D2�~ܠhmf��FXà��_����_�v�nve<!��447�PbhR��3^j���_���<���et�~��3Q���a�4��X'2[�ǁ��M�w!��2/.����}�Y�{̱��4|V~�n�..��21�%I+<4�ǰ��qIVZ)�bl�.���k�Ɨz;'=L/��"Å.J�*�k�@��hl����y1"L:�w@���:�5R�okcfW���@3^c4�	E��l������]���5�"�3$�i)s~�3�~K 9|W�4$���X�3�@���lap�q`�V�s�_֍��v�{:�H�b��}n����� *��{�3eúx��ދ��`<F�c</���c�,g�L��}kQ�5/<L�2/Ϙ��+%3H�E��펶�DO�P?����;9�(��GrI���b:w���t'Ŧ��)YFզ�;��ħ]�
f�����Zx<Z�ݠ	�\��g�U� `9N�O���G�"����:"bO��6�/8�g$��Y���9�rx��	�?I"�WTw��*\O�tc'��1�
���Ca����mO��0 ��X.�]o�5�tM�l�m�>�5�壘���yrh�^�'t>�lJت��iHh���Bl�|��Tu��!V�V\Ź ����`�Ƿ!�?�G0���U�|m���w~ol����)Q\���D�C��*�p)��z��x�_���h��g��;`�\; �:���|{�/n�m��ln@g_JR�ټ���P65� Ob�(��'yRZ5�#�` ُi�H�f�_gn����2R<�pV�,1���w��k�,A�
&��ͱ��_ঐ�ϒ�����գ�	"�;Z���<�0sX���{�>�Y��s��5�O�`�(`�-?C����-k��2*��>$�3�9)��{��=*��P�߄�1[N��6��
W����U:Y@�m�?1��tn>��ʗ���c��W�%�"j0n^<{[6�HTz$=�g��
��d����D[ϜS��D�+<F��1���;���^��ʐmQ~[zLG��H���cR�nr-m�Fb%XJ�f&�/��&��y��:��*	O|L#�\x�3������=�k���b�����{�Y]W�-����o�˲����o�\�W�1�s�l���d�t�K�w� �n�_����0�]�6Ή�XV�?�|r�5��9~6�
5!�H�78�kQ�c[Sa����4��ě��3Q�O��#M�u���)�:�]�����(��~;s���"��	șx�x�O��Za��g��z�7C�_٘�����n��3�>�tW�y�J6~LA˃
���X�^�+a!�Osy�7i�Ծ��	*�|�@f@'B��(p�E��@3I���a#\��ƾ�/�-!���P�M��X��a+�n�T�z���#HX���?�����+�n)_�|U�m�}���8�7�fS���<a9l�DN�=���X@Q�[#י������2FN2�!�Q���;��gں�����G�>`;��l�q�ot[���0Q��칋��*I���4�ˊ�֑k�)�����)�ز��9�M��iz��֏�:�B�=�#u��~��[5�a��,�t״͵�`"%��P1[����b���q��t����0_�\�uɌ7��=����)x�����Js�f5���r��g�����$�F�
P���<7�ET♌@K�	�_H�8�] �M+~]t���B��՚�i�iGfe �r6���R�����j3�A�;J�4�3;�Ho�6����Ry���YlCó9˞��}i��"C<��@�m֍�'CTGT�7t��&�{�4ˬ�%� "Fc� {ʹb��3'
�w��8ƹ�& �����-/N���{�M*e+J+��g54���GX��ݻ,��$���{��YA,2��m����X����	0Wl��;:�D��|:y�ÎRǕ��h�P��	o"^n�2uI屹[���v�1��d��-ð��!��l����#"+)���ՔI"�O`w��'N�����$q�,Ĉ��'�X2���v��+9R�n�G}V�����;ܹ��V��q�ߊ�g�oFa��^�����A����"��
�ٔ���C嗉�t�+7lV���1Y6=KQ�2�в��������`����h3����?�p���}��+ޯ��V� 4hDI���K]-!YW�' �Z������uFm�C]��QyⲌ��[���Ʌ��Io+�R`0zI�!�?}>�es�"DC:Q��s�wFʬ�%b-��xv������+kX��r����Ь���o�"��!B!��]	�{�����>� " ���� �PŇ�����)=)�7=�·�)���,eb&4�Z{��-\S�w���i�#�F��¢n�0��[�<�qK��}WZ�r�cdM�:�Alv?�>��aT�$��X9=!��u]:�[�����.�^�4KL�U/�1��*�����yՄ��@�3	k��ǌ�l�[��-� ��X&��T	Tݡ�B�h%�_�D��o�v��*A7S@-�ِ7�X� ���%�����G"�2��y��/w���ǓB�)@�\-+6DcU����EŎ��&`Oy�꘰��tZ�%a�e��6�5c'A�kYa��� ��b�y��}�A� Z�} ������*.��<r�K��,��|��'�6^�H�J:�<���aS���1٫ֈM��Wݵ���Z~q��Ѓ ��+��>S�1d�P:��U�S��1�#����C�� -�:bA��$��L!i����$=2U��O�����[��tt��[��@m:b�B[�є���7=s�B�l{(�f�2���ު����9x_)�e�K�bG�yo��^�������@,�x�Qi��rҞ�{^���� �]+�`Nyy��oqrJ&K�X>'�2p���k��Wh�T��F
1���E"뛣�gP0�\>	������4�$�ƺ�9���%��~�6-{n�pE%r�I��|
����$���Y�t�3c��WL�H���_�-�l)������=LȻ	J�K�,�������S�rw�F3���L����SC��i<Bh�Η�֦V7A6�q��u�Q<�x5��z{2 ��ꅹa��r���?���y�A��V\��q��g8~���빃����,����=���
|����v<����G�\#�-���R�o��j��Q���^%�Z���#����
�� Һ��4bh��(���W�/T�vCf���pK$�e��X�^�� ao@��\��6�b�_D??˿Q9'�$�e�7AxO���;��/ۊ]a'g"FXr�g��A� ��Z,�/c3G Yߡ���Vou��G}=����Cve@q��֮���&I�?�5�L|ײ&�6GۊʈKO0r7Z�X[H� �)9��6nn�@Tǐ@f��!9a�V4�ҍ�H��͸*�fq-�{Ϋ�(wE_<��~�L��>n�_��e�/[����z��3�����c�4���|쓗��>�W�7D|_0�Ґ/�d��Ѩ^�y�{�Ю��(-�K�`�Q��7k���ªl�2+�/a)ݩb�t=�V�ƈ����J���"���������Idh��?�%�F �)m�d���B`ftLd�'�]w�>Xax7k[K"ѕ�$��9����j��3��p���2�l��<
GVzvOP�vʐ��k��k��v��~�#�RW��A�X3,|X���(�}M���E�Q��J��ͤ^�#�j=�yg�����i�M�8
L��c�Fl0���-LڭH��>=�eG׆޾ź�F�Y�K�YX�Uu0s�ѩe�"�	��S�nt~�o�l�mgI�X�_k4j��(:�Ɯ��{�P���oJڽU�5�̑�	��^��]�ŎV7�ZT��S���r��Lf�	T?vr��w�7�eE!�y҂Lcb7"Tþ���
W=�/&��g�QZ�����N�/St��!˥��!clL�+?�/��65ۛ�
�F;b+�)�k�Q̖�z �o�k1�F�"��Ĭ-ъ73WC�BI6=4�6�I�A���rk�i1^s��HN���v����� /�9|3a�o�t�0ؙ�#iz�BpH�#T�Sc�y4�0J�����+��P�iL�|��wSm���ľF����J����N�RR��n� �⻟���T�!��!$�+*(�ӡ3��,�σ;ֶ��*��kI�맱L�Q��\���2X�9?�@�^<:�׫i
��t/FG=���{��oy�y�˥�10ޥI'������[7>a��m�>OW���P�ІΤ8��yQ9I ���3X�Q�;��� 7�^��:Nn'��&�{��7�V��F^>�q'���ƕ�̥�>��W0�����~��˵:^4W�7�kL	����D�`��B���+?H��6|�'�x��L��x��m6ӕ=B�X��������oU�(c���ʯ�c�$ۉn�|�d���:\�E��f��G�]��wm��2��d����\���1:A��k�cU�-򣁕����ް��>?�Q �W6�5�1L>�?Y0��v�G`�ٝ�wn#
��-���?��f���v��O#b{�t
�F�C�]X���O�X�/���T3=B~u������PøRY��Sl3����Pd���L����U�Vj�����p��kr +�9����/�.	� ��RI�H�B)�}�y�4��m�rsi���gM�ٹ����g�F#����G�=f�s�8��A���Ǟ�D�rR�=�>;�5'��7��d!�/\Jg�'�M�w��tzl�`�b�EQBF{�j��ř����r&McQ���B��Q�����}�B�X���&ñW�<\g ���3?���=�w���"�/Λg�z?�= G�)�!:�^rV�#��g�C~����@6����G� �<��ZZ�HTT��h�OH�.��<���.STH��tZf&��le�l�gh�p�y�(I���ʏnB�j&Ϸc�ȁ́yx.a�۠�Q�Wh ~_m@���ǉK!1�_����$��չ3l'@�ɣؾ�|p��̶�K��LʢrA)M�����4߯R�-B��Fot��VZQ�|e-�׫w��s6�=��u� ��8W��+\��%r��*�C�sĤ^:� <��=��9Y�͠GV3�^��vv,��,�`�&v�~_���V�ܒ	U�d�F��V*�oca.QGG`2#���
���:G�[�憭��L��B����q����� $��GI�s]H�1���D���y�n{��t����(hQ��N���x�B�Ҟ�\�
�XW�*g�7��/EJF��>N(B�������;���{�G�9��d�q�hF0��#J��X�Ø���!4��W������4$��Q�h�8ٷ�I��f#j_�P�C��ÌF��U��g����.�!��吋Z3��+���%��S�Z
VV#m<��c8�`���}���Pĝ��$͈
]m��-J����7��&�D)6\d�u�K�,_�VK�lh�5��I�G��G�M���/���j�S�Z�'��0�k�Q����$�� ��o�o?v�\sƄ�7�amR����խ6%��2�J�r��FmB$��3"q3%_v83MM�B�g'�`�Vp�)O>��K`�pO�[�}v�{|�O��ݏ⣒��"	%M<V��>*��]y 	ŗ#��]d?s�ҝ=<�a$琣������eѡ�8Zi�����G��:��М.W܀[�\���π��Kw��b�={��O�1%�T��4;U	]��"�|�uDϖ��o<E�S����-�R
#�����D'-��������V��-z���]�ۊ�=^%
��g|����. ں�tT�M��e:���/ӵ��yz� ZxW��I�җ����.)�G����Li׬���@���P������-��/w8��v��4&�	� ��������j%6լ�e�6k�����>�m��~�����RHn	֥�m�w2'XE
��ֿL�Ejc�َ��	A�Wr�oʟ�t}�ƀڣZ,����E}�[l�g��.'{ܶ^$���{�<�Z3�q>�N6��x�C�@en��;g!�[�;9�P�$�*�bn/hg��q���Ϝ�{��Z|�_��q�u�Q�j���Y�=6�cZ(44GF0�������Dl�Kڋ[��G_w�EW�?���A�Y½���(�4�.��TC��¦Yj������	lNu6���w��S��T�%�,Q��A�bd^�* �e��	� ����'չOe]%\��Θ�O��)�Sptl�%zaX;�/c��J�8L�&�d�z@<jԵ���g�	-�������;ߨfO����0��r}����bzJt2�'�V���=
�.�P�9t�4al�Z��(Ґ�U�E �ݖBYZ�ܺ�lMwҌ
��x��ջt ���g�*:
�z"�������ܛyS���k��܁�`8�^��9�y��ɤoE�a��6R�1�{cήQ���-	td|d�	����Rq��!҉ϼ{�'����*���0'�!RP I�)�Ks��%�>�C�x�UG�꓌>���w�m�8����\�ia����):X:zR�>�/��y]˗m�ӌ��ّ[�*g�]��:�V����x2X������~�-3$q	8i�y^#ʀ~����2gH_�bF��=����,aF��w䩭�����,>��x��jg_������(2��xV�ϲ\l�@�\-Y�J-SIh?7�\ WFn	�]��?oH�!>f�/���3�Bs �������.�=«�l����׎QIB<�.��H���V"j�k4P��0jK'��ӭr󏨜�D8�I��,��x+0gY���s C�b:�2�2���u���h�����pq$��h.;X���?P2�;��R΂����3(�
�|�^-
$1o�/�/1�t��tH�}���%^�������/7/Dh���,�qBXs1
�;
���]�������$�b�	��ŗ7�`5���.S��!k[��E���σH�x[�����6S������L��7	��v���$mrGIǮ��8ѯ�{���}H[l���G���U��~�,.�m=NdP�K��ռY�?T�����!�}h�Nc���6V�rt�:p:���i�;1��P�ϹY#x+���sĶe�W#��k�Ed3q1���74���]U1l����z�F��t����i�h��gg��k�m�ϙ��LH��^�����a��?^6/K:x�̈M6��gZ{:��ǥ'_ޔ2�Oi�C]i?��lO<^�F�	����j[{���B)մn����?�h��K���5@u���J��C?�,��]�����:�9k~��-K\3yK�{��e蚬�'�L 1|��� ��)@Whz,��'�i�gL G���1@�	��)����*ޑ鉰�f��J��w�,�d�Ĳ�.���$X�o�\���Q����J��S�ߣ_�(�G�����^l�����Xۋ�
8�zض�����2�����/�8?!��TRb�o�H��V?�P�}Q4^�P<#p��q��ĉ�oy�$X�an��* ?���n��[�,o+�2�7F���;y �l}��I-�V�ȵ��{. ����l��H=�9,�;TC�jS��(-�}8$"$������(a�����I8#v�\�،Qn�V
�x	/d����1�1^do�9��d�i׶^SZWS�i#��A #�i��F��/2U���}�3�ޣ��N�+g�{�"�	���G�	��
�h����޷P��?A�K�����诂E~Z ߱�f.�~\~�;�e��>�-B�Z�G�����u�ưC^��X&i��V��L�+���)������(ū� ���>h������`�Q�ALm���P�)?{Uի����w3������J�z(�m��8&�B�͆�E=[8�_s}���+;Ȧ�٨�zQ/���UX<eT���.~wF4n��dy�nn�*�l��k��2��o�*4r�`��uo�*�"�_�����N�s���q����oy���sr�O�u.�׿�o��.ר���0��=t_j��;A_`�~�t������As�J��8��JgU:��W�v��5drj�e� ��+������zK�E��Vv��������<v�ǰ�c�7����	�s�_��R�l`p�W)��a�{j�UGUHaD�/I�iAbQ&���bku�il�L�^]<�M�:��7i>��ܼ.�]�v�}�L�պ��ۉ��t��F8tJ~J�z�V��h��6b�̪l�F\�d�t{���V,:e���x�����T�1	��ȉ[�b�m�f#����h�On���\�#�v��t�b�r�lQ������	��`ث^�!�vQ>>-���	�66PS���6���Ц���Q�P"�i
)��p	�hxa ��Ғө��u��%O��$����݃N�7�6����)g䏺�^`V�D�L$�bc��
�~�A/�:�,~�Ҕj��o��Y�<]0���$�j�&Z�o�9��YK(�0/`?�8P�~M;	���wyJ����n�述q �&��NNՖ�K��7X�.*���rپ���"��`�5Eh^�P��4vc�9�r�����[�D}�^��X�y`^F�8D��J��u����y����X��zӗ^*�_z��_s�m@ƿ�BH�ԟ�EZ�|���Y]�����]$�_�t��[0�J��.��Ym��J��R���5C��YOMmkɈ��݊ڡ� a#�z��T������(}��*"��"��F~��4S/y?Y�9�b|l��~P3��82iI�gĭ��H�P���2̘\��]F`de���({� �aE�m������ե���%���@�p��ڶ���d)���ϋ���	�ԦX��m�7a��6���@�H���y_=���l�c�O�$��o[����F���6��a�̂��$K�d�<lI�aE���L�G���{�v�5N���aّu�����^�M&K�=�p��I�{y�w�9�E�d�@&�{si<'N(�ћﭞZ�nS��) ����[�-N����v��m�ʴ�Y��SDd�Y����l�Fʴ�l-ۋ#GD�*Vf�L2�"�C�;HX�BdZ�i��S}?��:���@#WX���5��Tʆ�G�F>�c��@�U�5��z�n`$ݨ="���6�%~��$]o��=-tlE��<5�s���<Ό�ɩ��X4�f���įT(�qM����-R��%�$#��jB��
8���G����LɈƊ�p�.�(��Gs't�T��z�1W��hOv����'�U|7a�{A֌��Ϫ� �Kj޺���r�ɹ���҇&�:� ��C��4���@���/&.�ol�H����_:X�|ʄ"-!��T�}q`��^������c���yr���(11���v_�4��X��/k��z$~�A<e�T�%�k�a>��^C���[��g|.�����9AK��H[�����'$���?�r�$�Z�?���S�`����S�G���CIA�D����{��t����hb?ڀ��V��V�Mr>�م��b�% ����L�G�Հ�D��	M�)[H�e(c�+O�Q�@T��wa�c��A�l@���m�^0���7�g�ps���)w�4nۀp���������u:�Et\}`���^�ׁ/$�[��c @37�YQ�e[�``���j�*�)膹L2u�|�[|U`͇r�-���ajs��H�q���T�BOf�?�tw<������ksUt�0Y�!�h9���l\魶u$�s>��������P��4�0QN�"ʫ�|�{J�x-
��l+����)�����1�G)p%	%�V���b蘭K�`#���F��;	�}���;��UUK2�or��	�g�r&���>�4Fot8��*��GY�:����L��ڶ����~���QK:q����D�t��:j��� 9�ȇ�jQ�����s�B[�� �kZ�.�W�a�;ykcWu�e�~/�X��RfJ�LW�ݾ�b�B����sHH��&rIn��	" �p��|��ak��v2�js� � Yg|�X��6o����Q�I%�c�N���M��E6)�u����[e��j��J7���q���|�� �F��ܺ���'�{���=^��wM�$��3��t����B�H���$����+*��g͆\;>��2��֓�)��硾U�g]�CdI\M��f�yd����z�|�$?��i����7���Y��N�m�m,pgm~J�|qt}ć_�d��j=)<����s��],hn�����v����b1�#�Ɉn)"&u�]�|*P�e@���5Z=ɘ���y`)�R��D6q�Xx_"?��ačq�2C��/`�6���Cy�>[�׹yEîxn}Փ�.����ڴe��4"k�-aB�?��+�<��6 +`�J�g�oVOTN/@�
?�	dƩ�$���9�-��P�m����p1�s����e�: -`Sh�yQ܇)�n�X;xK��iM�N��
V�b���HIN��&QS�@��!��� V]-�ݗΗ��=Q�{�;�SѧK� �N�Z��VengGO_�F�
��F�4���_�=�X8,�G�N/,�JbU3�c�W`A�X�35��"ᆑ~�����/;҅�m���>���`~��@QF-y�c��!C��]�s�+�Y�ԥ��F���fh�Sy�� �֗f����s���6� ��#��T��$W���i\`v�l�E�Ǆ8���yU�'��}~b_��c�6��*��ٷ���/�`�m�_���J�."fK�h����c�<)T˸��u=�W��_xű{��]�18Y�s9X\�y�/_����	D�����R����߈��e�G��±-rP#E�ټL����̷Z�GR��(��+�1H��EY�C�-�����4��S3\^qQ�������`K�`�A�L}b>���	4p!�9��?�⭬�u�b��S�4�y*�T��,s�G�w�!�飴�Q��t1�Z��L�`�0f�2�g���]C#Sg9p��ͺ�AM.zi�{��T����W�>��؎��<E/��X�K�D�Fy�&y��Y��ѩ�Z+W&.E�V�߱0�g?�p��T^^�3$��"�	'�T|��X��o%��-�����`���.`�JR@RY���x璸�l�b���)��	���bǎ7�P:�B���7�h�LZ��B�L/��G��ie<��x��\v'����Mٙ%'�����b�n@7��XUt�a�tYU��Ϩ!6�#�����b�ҏ+����7qCȳx��:P�1�Kʂ��ҡ=S��3�=����Qd�(oX;NVҕ�15�F��`���y�IĂiI�`�ߏ4�:\�?~'3�����P��A=���ޙ�%���^¾w�0��x��C�������E�����fYo�_�<�o}"�{km���y��:	�J�������8sa�R���AU-�hJ� �7T�+�9��`�M\��Z�~����j��7�f�i��^jO��l��z�
a�k�~��7�1�_�[��E��7�{����#�ˣ���V=��f�E塹s;2�<U9zho�6ԋ��8�}X������������� �[:!���t Ŋf��#l�~Ƶ�vu@0��dR��-2T��=�O�M{��^�yX�gn
 �;ؙ�����:
��y�����)#��D��T�=��R�MK;E�s󹬼�I��D�bm����A�la�e��]]aux��q���d��Dhծ�ط��/�W��t�(mpl���Z��'���������S|E�R���Yw�QkPڴ{�y��e%+ǳ�L[\m����-�C��*��O�8,��'������"ĺn���`�+ۖ�1w�S�OI���g�����ud5?4�	�O�s�~��=ڎ*}S����e�
���qd��I(���*�f�_�;�6�0O�Hhk��(6�wqu�y�$ј��Ƭ�Q�v�����0CD�z4wA���;����T'Z1��E�X�0�[38��n
' ����J>���7ɣ(.n@��5)y-*Ǥ(�Y$R���������YOx����V)�bP�e�6�]l��LN�9#u����Z߰v�\�d����H	.pR8ԊC,U�ٹg'A�on��;�T��Mm����VR�T�6�C�]�A|h�ypCF��z?�#�6�$m�v�]��w�����`�dwٹ�cY�q�}���]��66��~ECL&�����/L�a�N��=�ĝm����eW��:��6iQ�fk���q���I:5�bX��v�#����߼/�	#7SM�V���������Se;+/�\�3����Qf��m�L�Ǐ��+�����o����
;U�%1'��+ �}��#��m=T�z�S7l�*c�K�R�e�ϋߑg�^s������P�*NQ�����A2�&�����ξ�cb����i�K�di=���C% ����ꥶu�6�o�7��G�����I�]�{K�F�J�U�NO��8�?u��k����1�-�Y�+φ�xl*A)")�i !�%���7�<��k/*�Ҷ���f�c6�8��bQ�B."�����G.t̸�/GnSs*�!lGvx��1e^��d�GN�b�Mg�l��p1��
T�-����.mc��Iʵ���~� 7�vy6��� ��ڭ�_D��~�ŭ�4��mi �mB�^�����pN,%ti��Y��$�V���
�"���?HTz�׭�c�[���Ԉv��0m�Aҏ�31J1ħ�V�f�X�B0h6�E��mec:m�,,��?@�8�3-Q�Ν�Y�`��u��d�Ap���dHfGP���/��k-�u��v@<�蹽���Q��d�l.b�g
;�W]:�����Q%��!���P�~$nE��f��'�߰���U"C=7��[mǃ�|�1�m_Bj}Y���!��S�4OK�u�G�cO��P��U��t7�x1�iG����"���aA���a�(�bE�}�����R��WG2�6⒮��H3+7HO�J�~���wX�;�@mT�ߌA��P�!1"�5!���q ����Ӣ)��ٛ �l1�עM��(����@bd��x�}�^�`�>jr�Ɵ�����!�VjP�'�s��a����NF��Ø�m��,X�l1���C��W>����Ħ������]k�����_2��	l���Ԯ**��G�tHY�u��L�5fi��eTl����v;3�)R!�eq��W�eZ��G���ȝJg�l���'R��S}�C��ֻO��ƒaqM�S��z�lj(����J��@V�#��?�8I��i��L�PM�i����R�@]x���A?Һ	N7��ִ���MK�����6S̙���a�����$�m��|��֝b�^�Z��g����Oل*g���� �>8��-]l5��oNI����CR�9�I��
�$o�,8��Ļ��l�`+�vWzTRuG4�(n])vE4�[893p>�I\�ݯA�����j���(_͚z��o�)��DQ��V�ܒ��4lvurD\.�,ˡ1��
 ���ɩ܃p���7�^u�g�q��X�Pu&34��� �O�����D�
W<��e$�����~+>-@
�X�<	� ����v(@t}`B}$�S��X�|(%����毆	��U���KG��5i:�(!��IY$[�av���#]�3�1Ԑ�őr�!xa�����6a4��∽A���\�����J�"(��2Q/>���,��9b����dB]��_$���}P"e|E铔ى�hJ5(uDY��7|�vGk����~$����DK\�,�p�mvoP4�#�?�3����)�#��5w�f�m��Ɍ�yCL��fx3�D�DfQ�y�jV+�W�cҘ@,*,�۬�S�ߞl�~����ݮ>�%�5�����
�v�s���X�)���ӆ��л=r�m���קqo�K��m>p%:Je*f����>GNA��e��C\+���줲�]�����%i���R*��C��M�o~�U-�����k��?odI�ũ�J��ÿ�K�x�D�c�ր�D���7� vG"Re�[���uW�y����r�4��PHZ�BO[���?�87��b� ^DhC�����_;�� 8	��?��?V*b�r��;]��.�N��Q�H�-.R@
9���Gx�%8=9`�3��sn�����+Q��g�G�����P"=�B�N,]4O7{�Q9}'�VW]fV$�<�o�fc}u�%*��=���k'0iN=�*�ҳ�������*b�H���w�-���c3��S�U��2��e�䔞�����\h�� VAPJB͖9�ޕ|sC�Sw?���+��e�!�4�"G�r�x�к�|ďO&7���V��-K�S�ie7�]�D���[��N> 1�L���� 9��Q-d#kˏ��%�۵KDҗV@��蕎��U�L��"\"]�{%���}'�$�aUǚ��5^�Q�6I�$�E#��8a?ZY��:��>S��zm�}:^�[u�:ᕰ��x�RN�n�S,���pL����fͽ�`�c ����*M�Ci1�ǆ�!�&?��H����%T�6%(��#18��xao����z#*�c����m�l�8�.P��Q�v���L�����r�$jm;T8����P'��)�-Tub��/~�k����r����!wb�ٓ�k{�EJuP�
@�j�r���<)�M��X�FU~�4��Z"����]z龮�0��b��8��N�Ϩ!޷*�
���[ek"����g����Z��v=wC�ɔ�$����S���٥�_k�H0ߋ��ƚu�&����K䀈�/a&o��ލ��������Rt�߀��M�����^ܙeX��\[��L��" H���eJ�o=��~��O�Al�l�
�4�sV�sC��(�ֺщf��*�j�c���9đ�� �4�����}�u�T�(EsHR	������P�z���{�m�����'�]�S�5=WӤ��l�c��R$���Z�|����D12��@)9�hH���Z�{�X�XE��
SYuARc�q"6�2]�FOoη�����`��p�B`��<*�1��2�#�QQ�Ԃ���O��-R����Ě�&���ݿ�����ο���7�Ȍ�dS�c�^P�� /�JF�=`���-`���7S�y�D�hʍ�ln��S}����8oLb(��ݽ,��lá�����NK��g�f<sĘ)u�lU���ӯ�.��.;q'~���[q>P<*��c{z��C�v�<t������v�6��$��~8�3
�t_�C��>t��2w%�C7�>�4q�ImOE�7����/!ʃynj�zZv��wpDe��?&%Uvc��(z�ܴ<i�K����M{�Zfr��P�}�vW���ߤ��lnbޔ�n:I�KH��.�3X4��9�h���&<�`P�K���u5�Va�W^���Y�N�[W�فP��11��>��gn��P"(QьZgb���b�N�k89(�xR��NP�m��m��R�?Te�qo�xb#�� ����M�@�_jH��ƊO�%;�7{c��S��~cXX3��<=ޒ���c����r�	�c.h��c��_~�4Xl�Uc^��߿ah�͔"��$^h�Y�� ��*����3�Z�@�1��<=��ERG��,��g�z`t3ߩZ��lP[b��|�^����Ԭ�����Ï�C���ڊn�o�n����9����(o�������:��g������=���l�

E�A,�怼�η颛�cۚ�s/��D�˻�rYeL�e�a�MQ혨۝aW޻/��?&��gQ��lWC�$���J�'���n7Et�2�C�7~����p+���A�^ۖF	���Ȝ� 1ZH�c
����Ʃ�	�@-�~�i?�T���%�B��G�d�D��xw'�J�j�&9�3(0���M�q�sZDV�w�~���B����/o�d��-v����eTT@\�]砾I�hX���i��`�ܟz�X
�B�~.��p�jDxq+�b�Ė���-*���ؒ���I�섖����a=���}L �&""�����6`���8P�A+���a�&a�~�'�HI�x�PE���w��lӸ��!�ɦG%l�SJ�J�/JH� s.��8��m��� zbO��[�|O�W8����C�xe���.$UQZ`a�4��ۣ�f����q|����2�ztb7��V��7z*AxH���I-�Ǵݩ`�dqߩ���dV�7Ů���o'���0�o�Tv�TMU��Q_���'D��*��g�������mHt�b�~Lr��"��느
"Q�4��ٸXHl͍�鸖��&�[��X�'��+$"�lY����b�I�jQ5lnՀ��ۗ��P>�ׅ���&�0���>w��oD�S0�+��X�?���tø���/ ��:qw��?G+M�J�K�����)pg8Q�N��� �Ty#�5�X��ǈdGa��/��0<�`�o�ħ�����4f0i�����G#�p-O� V��?�p��i�뱘�|x�oY\l�@6C�TQ����O�����?���3و�/��������Y��� 9�+֖���0[�ɡ���Z��B"�`���أYD��L����Q��#����YL����rq�
�Ii ���;#�S�H���y{�������!K�z}�J�X
�Ҙx▊
Hy _&��&"�����u���Vw�u7��B�&��B�+Y��Mh�^�/PP��G̓�����Y:+CA�n�%��֎�7�7��	\c�:�u*���M�2���o5��(i�!7�7EN�X���2 F�+���WKM�x��<^��'�O��SMw��"��M�kE9���4}|do	�/�'���@Q�\}]����[�;ൢl��.�6�Z(<>�J�.h'�=�ڹ�����������e�LK@��d��,�X����ALxꢹ���ߦKA�?�ˑ�� kť"b���W�;Z^T�P�{\zyÛxؼxEVe�ŔMF��t�x߲S]ۣt$�U��ư�C,����~���&���)��ӛ ���CDKФl��+O��POބ��X����
��4��퐰A����b��*��>�Q6���m�,D����͏
F<Kv����u�!���h+��;�n�}%���,DY���ޓ��)ze�d�O�]���$EW;\u��W���o���7�F$�8�<�`/(��E�-�Vj_�F��E��T�=��/���
�@Eѳ�-�|�v_*����2� �?�0�7 �![���0_��SG���$����A�K��j�`0p�e�@�t�YjS����}L��@�WϨ�N	�Iq�G�jd�]л��Љ��cw�kx��3� f�����Yu(y��(��ș�ĞW�)�{����_baWb��a�<(�VF_��^n��.�R�?O�3��%���?�rM	i��L��^�Q��)���
�w��>��'49(N9֖�<��W_=վ�"6��=t|��ޢ�Y��^�=��qH`ia��ngr���H �mE�P}��a ���Z���P-}�Tq���6��f��}9 %_ V*��8MpQC����$b�?z��4�+,������7$@U�y�H��%F�4�`p�$ŀеE��WWߐ ��Bx�.��$e�|���wF}�\�	m�3�_���9*F���U͹���B�.(^L5B���ODpQ1��bb��a�.�\j&S69�%�0M��y��3��^��
�}嵐i~x�{��=wP��Mp������Bw�c�u�����X�`�U�����M�g�4���#�X�$��w<��pȃ(�ٟ�����#5���@�4vm���L6���?��J#�����8���3��s�b.�d	�c]��렉َ��b��w�3n�3�`^�͑M!"��a2wo\~� �xM!���r�A�)���U�HjC��}�l�G��M)�ƴa��HC��*ۻ}*�[��=��%c��]���uw�����"��B[A ��*����I��)-���w��K{TWIy�w 5�+�%[�7��L��2�Ɵ��v�i��4��X�/o�yA���`�]��D�}Q:|�u�z��ꂌM���p+�H�|��L���m�]+���<�=N��y�w]9��qv��j71=�V��OgT�O"��6�Rݥf���O"�k�xZ)g��E�up/U5E�ȳ,��QV��M����y��6\a�H�*�z��t ��3����m����18����(<YQ�ʭ�S�N�Ý���AF���<؞���%2>�n�;�s}��dQ�6��-�-�C�B�1ԸQ-]�\5���	
��� �	�+y��fU��( �v��U�����&t���p텗���}�'���ɮ�-7��w� 1*ecb���/mE�en������U+���z�XPq�5,6�Wr p~#HW�tP�B0�k9��*W*9Z9� ��9��o�=2��h�{&�T��5�ћ�t�)(%`��5xCY�R��r�ȦG�b��&˂�y�LT3�d����=��u����+�"�cm(����E��j���K�G����~gZ6m �5u�C��V�.���s��G���p3A���c�-.���y!@E�a�I
�����g-�d�����za��C�G���}���(�w��CCR�0cgj[E��T��i�Q�n�}S-a���1��(N��e��X��%X�|���w`�|M�w5n�Q��2������˺�%�8�k/���(�L_PM�4���Q�:u���%�*��Z�hȽZ���Ĩ��b�h%x--��6�6�'r�D�����'��Z�8:hR�՘y�*��AQZT]yT��@P��쪸�h4h�����6L��y�$#�Ar93���ѡ�ې�N�o����n�A��.���zMf	�O
=�Uof�~�B$@dK�S�W�s�$��Sx~RQ+oW���κ���pWw�F5��I���8G���Γ7����P:�_�Ĳ�5��?�w��<�`�v��lN�ڌ�N���-|�� %�.Y�o�^L=2��tT��a�w� ���[o�CɌ���e�B�-����:�ɷ�y�mX����	�Wti��%t	����s!!@'�*�q'F��< Z��lj(� �:�ق���F� ���h��ĜhxJ3��4�XZ�@|і@�?��"�mz����˱&���rxj��ҦE����$�N�H_Ӳc�pkt5V�{?C~�mqeV|��?�ѯٌR�xy�T���fld7���T2$|8�k�mt�,7���sc�S��l?qy����������rE{�WF!!�w8�9������T<��'�	?�k�{��鞩G)?A�f���5%6�^#xb�f{���Wؑ$a��kV�	�纈i�����~�����%��|�h��~抽�e����iT=$���2ǣ���vl=uȾd�4�����BVDN�vP/�-�'���\���Tόfh��Ud�}����	����d�>��!����n�l`��Iu��|�����#���e��W�!5���t��3�x�ӳ8Q�@���2�Boy�\�|�27FU')��Dp�,?��`��J4W�7���4������>��N����ۂ���ΈA���6Z�o"!j��3e��E'�	Gp������0�/0G( T�ڇ��hs�	�<��41��Ir�ֵtz�(+99���j�> ���
0Ue�	ӹ��FP�^r,� �u*YvO2�	a���v��K��n�o�I+��?�>�~�o��0[r�I 3@����I�]�*Nݒc�*x�,�|�m�G�#Nh<��R�� q
�e�W�2�j�9�e�QO��e��D&'��0�0�.g�6�+z71 ��o}����,O�ruĽHQ�õ�O3S"�~����&T���f_�lI
̴4��bEB���0Cc��oҥ3��i��oAN�P8G̷6j	�_vB?���>�Ƶ�<�EP)w	O�A��zAh��OO�J��x���4d�P�&kX6�nN)�y��}菞�"�Ј&k���6֏�����A��!�*n��V��Pjn/���m5�ç��D�e�o`��z�Ŋ�R�������@9����O5��i���a��zڲ-Ř���M��e��a�q�4w����3�%(x��V�7��^��ʕ�`��	�J"^@,E�/^rT�@�~�qF�P�g�"�?C������V�s s��H�ؼ�B��/�*��[�8&h h�5G���317�/���Z�9B�Y����2m�b%�baF�w�S'-ǚ�9f�9}s�iJ�@":�L
��/�u�ߦؗ���I�B¡+��}�Xmվ\۽�����M]'�7i`~�뷛�W>��_�a�)�\�V��D�%=*)��6��۽�͎oL"�~��*c;��b��l:><�nwT�L�D�YwPk�;���$����|����=�')�V~���նL(ȁ=.UDknⱆR {�4z���D�-�R-�I?�U��̫�i���Ց�c'q�E��<IPGا� wǄZ�-��A�&9�>d6dV��4K�A{k��x�F���`����xb�jA�4	(솋cx�K9�
n |7J@����7���i����{!����(� ���f
��[,"�í��T�r�[k/��u�=w_����|V����V��0M{C���Ty)��?:�45K�Ӱ���lݡL	�%���sI��	;�f���� R{Z�ti�c���/����ף�_�?@�ӵ�+������*�`$�a�A�<]����Q�%�����U��ǚPM!EϾ�����=/eE��g���фU�_'�)�������|.���u��S4��bF|��1Ѻ�*���lL�{>���A�Dm�
f��4&U�ԌVQ��k��;g�OMLF^�v��'���X8.��������,"P6���4�F������������+/1�O1���|�Mtq� ��G��D���89�S t��G��v�	&�_񨄶�h�,��%��������ޥ���j�U�v�;�/�q�ҹ��7pg�@S;�4��cv���!��ɬ��:yOnA��g�0��}�D��_lh�x���rX��L؈2��k�;�%$�+���[��0��L����U��~��1� �)"�e���zmm�&�To_��&���Cw4j���?�Ѐ���2ʍ�х7��QN�]�\]��̱�^���9��hM�0EK�E��	����1�}��z�!ױ��]9~S܆.v�a�����ب�p���q�������Z^4E�E%.�������kx���Kʄ���*C����x���łvT�AM����z�tO ���p�/�rGJ�0�5�x�|��,a������;T%�ԛ��:�������Vw�ƈ�Y�t�g�xp:�/=���	@)%�"�:n�[[��5�Q��ni<��T}���d�� ���� �Ż�<%;��o��T��d���@�ڰQF�,5����5k��5�C��,�}�H�-B�O2tr���9L�ձ>�vq���ך������/�}h��Iv�����Z����78�i%蓚ݱ ]m��H,��=�L��FՃd�
R30�"��͵��R�uH~��ř�.�&�t����{�����^"D���n�}+��������W����|6%,݅��*�e���`\�.5�Nu���ILt�מvկ�.�r������a!�*����c�8T�d@�a�SA'�d�������N����b{E��v*I�Eӻ����U���h��{-�0�'��G�t������M��7��Ӹ��mՇ��d�b��OBN��"uGעW"�O��ߪ�^���/��*@ЭZ{��:"�C�\���#O8���W[����P'���k�3�B��f��sTW�6��
h��G3����~�]�x%0�hjF�&<�٥&�f�wj�NB偳G`g����S��7��F��OF*���$�GQ����,g��Ex..$y��p��)U�L��fkG��(��de�X�\;�x�+t�+�q�3�@���J��,�v`Q�* �����C�fY0��W�Wd�$������:m'7$��q�BH?�D�bX]����h-��A�qPh��j�vZM�YY�Ra�;�ȷ��1ܹg�!��Φr�o=�'3�p�Ш���u��>��d���]��nH@5k�?�&�U�"����Z���)����YB�A��7���{s������mq��C�����rX�LG��v6|��:�Y�l2����
�O��^�Bi��cC�Ab��5>m��^9����wt��ѡD����!a=R�q?#�$+Pp��ZVĊ��l?u��ӎ��;������;aJ�0���R��°n"H�2������_ϬE����{��8�8�bXS��d�i-���Bǋ���'1m:�#|`t�����[���o"�/;�R^�_�p�·CQSk��m2��5� �F��ɻ29�����u�P�eҺ�Q�x�J�7Q�H��SFP�Ju�� �����y�E�%܀>�>�9�)�M��:����3mF��NWb{�M�F��(T�5��[�\4���u����d��r�
B�Ej[�~�8��^כ�O�qM�g��B��>�z��W>3}�^�U���ptJǩV���gT�urm@k ��*H��ˏW� >��㙶��e�ւs �?5���HK:��e�QR��+���_<�+8�5�],(��|#ʔ"L��yZ-���hP�S��8�rqi�\�H��Kc���Y�翸�����;�����p�a@/&�ƞqp��/�-Л�۪��h����a� R��+�Y�f;�4&�^�c����bs<Vg��4�1�\�ha�x��Ro(�H<�&A��;5���:i�hǫ�>�9F<�E�w���0�3(I?�^O�Th�������_K/T���S�6U��6��8'�z>W�_��ߵ?����^l����$}]�x�q��E�@����%�ZUo#rh������ڕF&FǙi�Fs���ҫ��@���[z�ϑ����힚���߲�C��)���$e� B��r�Zd�Y/�U[aY��El48��!�l���Ka X��������?��� 
Y���(�G]��&�J� ���ljF����AH/_ݣ_���}`�6����Ko	�����?�9����E�*$�A>c�eQ'
Q��'�e�h����c�~��h]�pg�u�D�ĭؤ�6�Z���p��!����55*�ūO����n1
��AXI]�#@��yâ���H�㡣�#�$�0W2qCvG�+$�.D��+G��&Lt+d�JC���;;Wj�?a�u�=[#,�rp��O�O3%������";Ԍ���]�]ӏC�� �֙}{U+��A�P���g��m#ڿp��	%"�q)a�}lE�����(-�8B1vO{.����\���~в���S^�J�
�Zu�!�N�9�:B�� ���P+t��1{�! ���g���c�色��봪�z��q���[��c+a�8G����^�a:�f)^xH��<��z�q��勜]�h�ܝ���]1_�qZI%Gy�C���]�;d��I�f��>�xi��h����A )xc���x|��.s��#bL�=���g�9܍��� 3�G9d0���A��y�| ���Ά��q�.a�z]|��<� ���z���K(�4��]`#�2�����h�gS��Nf܋s�a��ѭ =�H��2���Lpz�J��oa���v��/�<�\@�!�at�N�Ր/h�OA}�xAw���Q
{ŝ��?H�x�WbE�Q�wӗѬ�A2��3��j`�[&�<}\�]o'[���. g�>a-N��٥J2���S�űtD]:��)���:]���3���/r�U5:0�K�������'�C��fܑT0鋷E\!��z+�������T�~⭙�5 ���/=5�(U���5�x����"�_s.�(��:g��]�,[S[�s���q�<?��8a��{�%�2�Y�ũ�e)ۉT�v���e�!�@��ĭZ'�~J�P���vn�-���!����WS���(���S$��:J`ED� �����9,:K���cM��L@ &7�Щr�	01t�s!�Ɇ�)���t�#5�G�<�8?�_BÀe��k	EU���i8L�d��D��� �}iz`G��9nڞ�Nb��`E�AC�y���G���r�G�Қ-�m�y*E�
�_Q�,:2G� t&������\�y	��8��Z]�1�-�K0�=�\_P�G��`h4�>�Fh���$�{���A�ɤ6*^�@?x�$wm�Q��w�0�E�l���q�dނ���1/�ڲ�����g��\1s�7��n�=8[�G��T�DR�3� GQذV��'��f����YJ��΁���p�m8p��EHK�}XG*�d(#��
>�Qf��|ΪmO���y5o�����h�0�p0���*z
JT�(~�M����Z�ҡ^5w��}LvZ	�7J�@���4��lC�B���|m�gM'VUrf΅�e��֌aA�W�%@� v}(������=�bC�/w>@�1&ґ3������ ���^�o��^č�C����]����>u�fX_�3�s��aP�a��b�̨r2�`�&��|���?� [�J��Z�jp�i�qq
�\%�i_��q�
8�QgЄ�g.e?�̟K��
6��[V��S���^9�,���Dms����;�aUb�w��}2wm� T��rTC\�0�BE�@�����c����&jB络C�Ě�՗��il�hPc�*��4ʴKR�T��j�P�_�ߝ#���؊i#7�[�wU��Gƚ�	�K�0j�3�)�w��7{ʖ�|��E-�OE��mԮ�'
�+�b#W��
�t*�g�9C7@���$o�����1��K@��'>!��jG4۩(�����_c�N�3A��K�ɷ$G�N0L�����)�9v����jL�F"�e�ttϠ.7����5�
����0��qף����6�$��0�m�:�-�~;�FԸɕ#�J�����GI�u:�+�Gt�U�n�>}R�׺U6֑��j>\��R7���� �[���t�V�nur'����j�{AF]*�Ҋ��/�{�w�)��!n�įs��fmCR��K�I0AVEk���sJ�J��)f�����̈́(�	�	�wX����\�P�aax��~X�"߀P�.1^BH�t[��������s|7Č��Ƨ	�Z{��)��e���y�4S䒹6��`�?
S��H����J��;��:�9�'��#��b	�+���:'^�+�yg�[�)"҅`tU�U�~vĂߜ�ˉC��q�(��w�����RpC��Y�|���'t���U��X"�=*�;z�����=�������i5���Q]d��tl�!��t���"�t�^�l��%����"9f�}�fԽ+�_ˈ��Ї�F�h��8%�������>�n��L{�t�+وչΒŶ9�s3��05�X��Ϟ>�"�|��׈i�Ij	�r(p"dsC;��V���.��Ӄ�9�'���Oe�Z�X�$�~%'ˁm���	����z�f<�͊�\^8��}�CA�.��{[$?RH�'R��sBL�Dԥӥs�^Pmڢr��3������{�J��Qp��ן�$}�斟WԌ�{�*)�'���5�@G���V�/9a)�s6E����Fh�pL͗��;�����
Y�m08��hP���.�)CX���d�(Ht��	6Ulb7��o��M�����Ib#=����Cy�!�����qx����1����S��+ Y�@�P��0� /�m��W�倬���Z8�Y�]�z+���esQ�l$����@l0H�	
�n�� ���OQe=ϒr�`��폽�;��y�<��_V�����W�X�|7+*%���O�����]zM�k�S�C�ɤ����rF���+b��Z�TQ�M��b�-4�k�i�pk�s�Li�������k����f���ֲ ���o�t8G�[�:����p���Ȟ�XKޅ!B�c&zz��|�USm���>���=_2<���	
2&��QCT)}Xp�~����4�p�ƪ���+�M��������!�0�>��R�<Af��:��ÝtZ�/�Y�C/+����/��M���c
�
��~�إc&���d����:��#g�[+��^f��g�.�n�������!��(����R���_��@V�ɏ�_WeW���v�$�!SB��/�T�īA��!:U6ܝ����#Kn�*�
[��>��d���%���8m�#����W�>�����$ow`C^j���V��ӓ/5l�/�(Ɗ1���L���e��T�Q ��t����΢��VB�׬�c�uS�U7K��C&��VX��N%ཞ��ےd#���7nF�N��->����7�ᖏ�pW��Њ���\����6�	���m���f!�?��&;x�L�:X�lr����I\��$ ��T@�!e<9�������3�G3���.^LC�Z���rqr�=c�����c��P��W8��>@�����C��U���-�um����)qq���"B0��w:G��)l�xsS�A�?ǿ�6���)0n%#ȼ[M�5ogh���wXzw��c�?DӦ��M�6i�q�=*�R;e���O}���h,���/���
�5�vs�/�h0�Q�%������2!��3!��8�Y�̵m�O��'�4��8��A�u�I<�+��j�zm�GB���@/5��;-u�ޒ����i� ����(�^HȔV������Șh:�;f�HFr�$�#<�3,fb�����O��̍�\${~<��B�� �-��C�ݟν��cz�a�c�g�xD(߇�φ���&1��M��XW�(eo�&r�N���<i.�Z���L��b��b�7=�8�%Y��͇���&�W%,��U��n�v��~$�!/�Qt��دK�N�i��m��ZKp�nL�<R�ߵ�I<"HA�d�����W`d��9�HW���n�?�������$|,�&�~t	+����<�����^�RS������߀�t
]�l�'��<�xՔ��ߣ��Tșg5�e��pC�Dʑ��V�jQ�P��4�i��{:���9{��}3a�^�Nr$�����Y.�Wq9��2�O�F�V26���]M � Z�\��5�Ma�A��JJR�[$���~����<77�n�.�3�F��.�v�k9��ƣwZ%�޳��t�xچy=	G�����'L�}�� >ҳ���.;Č�Z���\ ��.5����w�8��L�2�][1w7�e��rդ.Vy�GiALqoO�*�͹�v�� �t 7��8Y�ī�#����U�9O�I��WZ�v��g����@��8��? 2)<E-vu��z&�&�>��G��*C�x��V̰�=�FtoA�OVw:v�|�ó
���ϘU��;����k�(=��{�\럺���r���}��[7bC�3��um��=��hdǓ.Т/�h����~ݪ�0F�ȩ݄겁��pǴ�����Patan�@�*b�}�K�b�Ԫ���'����j�됡�_7��
�����R��J�3�QM�^�h�z����g���Ix����2��Yާi��8���*������kX���SbqCL���r����i�]�R���OB�����qb`ٮ�����?7�K?��&����rȴ��<w�]D����X�t��)���A�̬�)t��[�Z���cŽ��QL6y����\O#p����hk%0E�`[�o3�8S� ���r���]K@!�̊��R��M���p'���/� 兖�8�3�7P(ݦ��8lq{_��f�i��)B��,w)L�9�0If9q�z)�XE��?<��z��(4=yW�sb�fW�{	��m�G�u ��N�$^4�Nr��,Ra0*����n�6Y9�פ��+���o�_��.��5Zq�,E��TP)~�\Ƶl�wA�\7a<{��
�#� 4���U{\d�g�OS={U.��N�����m�:?][|���D�h��	�ݏ"#��
[��7����?�ށ�i��)|�_x�����vT҄���@�9��T��&�zm���5���YU��B�o�m�����%����CM�$��&���.E*���J�M9�u�l \c�H)�L��䒨�N;���H`�1q~�S�,�k���LdK%��G[f�$7#\>A8�O��	(\ش��X&��*V׳����D����2���S�:�(�zt�3�|�Z��i�"��^; JTc0�a�!������H�?��s�̮��~�!o�X�n[�g Q]�S�l���5���Tu?��KO�x}�����B��ME��kH�vτ��⺳9~3pш'G�����Ma��y��{oT����^���鋖��;odf	�b9��x�cC@�#�?oN�Q+$����xM��ڌ!'�/���yQ�&4���'���__�������fhX�)���Btr���.�_���AHn�&W�$���g�}���tY�{y���}	���t�ے�G���fS��SK��Wv�7��d�gq��Y�����xx� Ȓ�����&f�r3
��CE���}����ɼ<�P��+�j��Z}6:F0������>����~�ߦ[2Tx�����y�ݽ~���C|a,o��&�~7���WB���ۂ|�Jے�#��3��cW���UCx*�{W})�i�J�d��Eg��������"0WJ��N����i�o�m�b�{��QZDk@�ʩ|�,�"E�N�x�����xO;[���jrU%��z���q{�ߒ��wp܁�I�-����q�������z�2��z��<p6,��	�J�����l��*�3�0��7_u��φ�;��f��(�OV]�v䃄$B�TT������\3t�M<ʙ��,\)���*"&�Iq�m˽�3�آ�n7?�W<(��(��ű��8��_؂�D�AI��Z]b���/h����Nf�q
]7��Y/�_��r1�+��Z�V�Q7�'u�z�U�]�H��^篲zh� ��4�:���m+c��q{[�`��	�)R��j�5	;j1?ଅV��j����'h5O�����4��z&�
xڥ䫂�H!
���ل�AL�����C�=��m~���r	�{��B֜}:��v�3oM�<p�� <�e7L�f�0
#��v���0,5C�A�c%t�f��	����֦|jFة�I��7\ē{b��-����*�IA]o��d��B���e��WG�ϑ���0C��
Tknx��R7^Ҩ�X���f���Ƚ	��Br0IB	@��x�w��8����N�ct���Hzר����|����zO
�u�ފb����}}�� "4�B�ee�s[�Zf?C�G��3X+;��lܜ� �=jQ�δws�o����IR�f2j�I�_��]�9�@�c�p��3$��,��<�!�䓀9w�Ai�+#ְŽ�f=v0�����<7��Ŕ~H�߇`(���b�uB|̌�?���^�S��		�Ϗ�솊��'zΛ�b5���Z������o!Qʵ�N���c̳����ʏt!����Y`9��i�D�J!�5� s!{+��r�;|1�6�X�/޴��W�6�c�]?w�G7�Է���Ԛ�"�|�C�̅�?��B�Y�H��J8V�*�o��T<��J�(i�Z,�	p^E���e��YG��i��*� ˴������.˝u�k�gH����/�3� �o!!�3�$�Z=E�ƃ� ����'PWq��Oe5�9J@��)o��ǁ�;�yu�l߻��l84�6ul���� 'rŁّ
�O���{HUqRL�ͨ�)��t3�P�fQ���2�)m/c��Ws{+G�W��R	��ʷ�Z�"V#0�sԝo�o�Bz;Δ{���
�+���=��V�fQ1���̑���i����OB��%�Y��(wdCV(�_m}�听B���a�]�NK��=}�O�Z<6L/�	�"��¨�$U���T�O���[� v�7˗�1��J�M.Ő�<F8�SHz����ךG0���fX����Y0h��kcP���sGn0k����˦l����^۾��Ѕ��N���)Pd�	��c��l7�@{��U(=�s�2
��V�R���(�!�br�� �Myk2P�HLhE��̽�̤4K��V�''_u��1�����m����!"աQ^��/98�KC`�~9n�yK�H��Az�}���'��t�4b��e^�����~�Nø[�~�Bn�KΣ��[���&-3����Q��<���7���'��Gt�ȡk�|�R��6��s��aQ�&�{|>�2���`4���'�Fl�ۯ�{�{��/п���}ͦ��]��18��X�H�ǷDė�9U"��P̻{Y�T�T/�b�k�4*Z��5��+.Su�<>2w|y��K1��,(���9J)��;�7��+%��ؤ���J8��_�}�� vYŚ a�)WY�uO�����k��F+W���\)H�1~�q�%��Y��F�3t��>���7!�x]�Ϋ��F���U?��1��&|�7j��SHUui�yv��M����'�!�M�#.ҡ��Ƈ#��T��jBh�_��ї��=9�n[��Y�ͥ4�(��qo���9��_��Bѫ�6���� ���X[M�o
�	�>~��~iu�M"|u�9��a*���['�!{%�$��b��S��(m��֨B�߁�b{�#������ [D�p��pD"�uo�5Ж�C(y�C��nGW6�\�o�O���¾֬Ͽ�&���L�	�����0���ܣs�V���D�M��9��;����&;�п��S��@T�*`y?O0LDf�Z�0����5�j��u+�nbrR�9k�P�M ��ْt��x����nvg��E8[8;�@���fLA�J�S���t�uȵ��T��n�}�������',�W�s?x�軖X�YT �M�|�h��u�:���0���[[���� ��Ŀ0���k�#�v$�,�C�W++P�1`s\(U'�U���O�����k�r������Kx���@�YdRr���!���M���BIB��0`��� v���ޘ�g�=/ i	��'��#o��6U���Zx��DIRu|�|�WkM:�Y�����.��H��=mYJꞷ`NK��,Z�n-�0k��f�p������䦱�����Q{�;��U�f�N	ss׍*4���Ca��؍��ơ=U�j����3������^�}�d��޳����2э��d��kR�K̎(o]��4�G��po���:�5Ʈ�����أ��L��"��O{����F��˗�}��vk�K�I�bpw*狅� w=��3��\��VI><œ9{�Y��YNՖ���C������@/F��2H䊎��j��o�$Q�1]=Y��*Y��@0�{`���D�F�fCC�b�٬ �Y�����O������o3<Sk���I
�9ݱr�������s�iA^	�/RW�ϨpA�Y��Ş!���i�F�:�^P�*��a[�S�|k���+���qo�V0�"J_d.��+�1T7�[/�n��8�{�fԵp�i�O�����_%d�$k޺T3�e�_kB"X-c����q�*8du;���Ks���K����;V�[��L_��r��[tB_�Z��x�Ã�Ź��4޼���j(�<����t�Wd��Tr�͘zy#��QB��]�����}�N�}�5a���O#�(�fk�k�)�%�+��֠(я+)�e������Y��b���������~���SU�<����I��ʏW�in5�eo5���/���0���D��u���)�'�f^�蹓v�T�e�*���$]�Zp����e�c�'�Ӝ�9q�x���M&YQ��D�B+����Վ�
���Y��W�����hIJ�i�GD��6Җ#���-!t圼��si���c���kke��{Qɥ�%X���ֳl8d-FWZ��p)�]�W`�h�٢%�%ť�Hw���}H��eu�����-��w���@�ʸoW�6��X�zs�O���z�o˻x�����H���_Z�g��My����:��r��l���hs��ĭ�K/�����?p��L���Fnˏ�.��|ւ1/���7yY�\��"o��|�S�3P[�&�r�gF��<@�k#��~����E�m����S�wG��.�l)R�\>{��|��,�C3k����ك4�v�ʓ�iiM�fT�a�u�2p���?cp^#Y4�Q���2�y��9�؝�#�.p�Z4v�eN%��~s���y)�B�)W��d
�R5�C��wI�?�&;~s�e�ȟi�1���� ���$vB����0�s���k� >9m��C$�������|OeD�3��6�j��蠝��m�8��< Ӊ]՛�����ʣD��y��:����?���[�F8߲��������:���P�w����+��(J��e�6oo�4oE�JS]���I��&8��i?K��:�o�A��s+�|�\:��j�ED�,
~��P`ӗV�Eb�<��~�����-�H�j9獤�\��K��i�/��I~{l�{q9.�Y�[���@�Ƽ��N�-b�$Wt��]���F XPK�x��	������ �Td����!�$&����v�9X{��
�U)��]�S�- /�9�y��p����e��Pח�VV���9�X�bWI��>��ԓQ�M��p�2��t�t�����bb59����n�0rS�%�⺌����9;�Έ�21�s9ك%|�5����i�-�+�< Ԡ#.z�S��Ff�S+�����	�-^\� �PT���ue_�Q�.����6� 3��w�I���
�|�uO�jF�PP��U���T5�x�WX,Q��g�`j@��M�*X}�Ϧ<m���%����3�2�ƪ-�+C��B�n�1�,3yH��>㠰V���#��eP�X����̏�>���`�\J�H���Q/*�Mb�hv��e�܈
�@�4���ӡ�e.��	�v��Q���[�B֎�1-�|(*��p�I�I5��D�?��qX�d�nƎ�,N�̊Y�C�����U��[�;
�VkZZ,@'�[��j����8�:`�H�a2����!N�E.�z����Y4��wĆ�h�j���R��-�	��"Q�K���1�C��������^�i����!�E���F'WTG���(��^�U���\N8w8��g��Đ)�B_����Ġ�B�é~6$�6vG��(=}��(�#�G �]�H]��̯耋]��og5S��=��t8���=z:.Դ�K�Iʙv�
t�	7PۺdDQ�:@�}�X�����e�c�2�*��������b3��r�d��}�o}�
��	�{�<� ����?��N	���*7P��K+�U��0���[ڊ�*�A]��ޘڍ|g/-^����-
 S0o{�u��o��
Cyyf.��1>_��rm8���"dV[�|d{���ԇ���a,Dɶ`8̪���׮�Q8�،y�1�>2~��QÖ�GL�*�N��®z��C>$]��d<Eyj�h����^i��ߊ��E_k�nN$��A~�H>�Z���M!�s����@�3��	*O�T�7�����-����Y�V�1	�8��`�m@����cv[êS��|�흋r���bX}�i��d_�c��A,c��8/�ܾF,H�k�uH=�F��e8��g���$�!]+RZ�9d���{�x5��- ��_1�/��Ef0���x�,ħ�m��v��;חٹ0����!ҿ�1U����	-$�y�=p'ȥ�C�y���A��,�z��
�t��0�v�*G0��9c�e����%�%!��&���we/�:f�8/�R�aq@�Pܩ�X��K���B x���-�ʜ��A  �m,���g���i(�lk�0�T�t+���S|�k�����k��
]�IV3�a..Q�Zsn�;�==�[h��L����V�1�z����/?��\.j5S�$3��^K�<5q�y	�^��A��-V��+�rE�H�<g"襕FX$]E�hlq�#�?@\*N	{�-�_���Z�[ ?P#�*��9�d#	N�>�^�N.+�c=-K�(B�������9'�D�"I-�q���Āv�ś��־wF �ٴ��6�_�z�(SN�[ɜ�^2����[��|Fr�䍇4�19ӥ-z�A�6s�f��n��G*��JP����D���	�X�ҟ��-���׼8�=8�uߕ7^��n��1���7����4���O��;1c:"P�W���nw�G��1|�ZU@�}cuX�F�Re�X��t����
)�[��� @�?�{/}��A���laUm�/<t0��mC��A@=����x�������`&�	���۠��$���)W������rX[����	�T�mtI�(��q��J?_\���X�9eʳЛ�{��B��MG��E� C���i��ҋ~j��/�桔ǟ�U����O�.���\Li}�~�o7"T��&k�$���8u;q�9�f�<N; 	��~�..X���C��n#w��P��oJOZ�L�\����2s2��"��|ʟ�=��,�.�>H�p��ymo���ߏg�Ȱ��h0����Qu7}���@��2P�� 3|��3���B�q8��KM b���H��6*���y|�cj+�4��������6�����M�Th��tb��>.Sb�cM���y�Ai壀c+��|�F�aQ�+rn?$v��Z�)D(ߩg���}�ۛ�y�On	NLY0W�Wa$da�^�?���Yx�`�1"B	�tY ����a�4nc�1 �V�H�M��wYZ�O;��ω>1.˜AZ���B�ܻ�\\Rb�S&aK_�&�:��6�/�삍����,!.����q�q/�[;��ӿ�(!����x{�--t���rm)�gգ�_����,\߳ˬɴ{~���s�8�LR��ٷ
�f���)|�`�5��(��C9iI��n����^a��J��>K*����/E/7���v���@�̱Hjy�K��(��ڡ�p����Upˈ-�3�n��xd1<v��P]��@E\"Oޛ-��w�"�G`�I
*�	]��Nm%
�/��H�դ�/��pJauR��p��A݂�˧�I���A�*o�:�1Rִ՝Sԍ]UQ�oR�3<$�}��ٍ>ͯ�Pͳ� �Ӈ�" S41>��\NE&��������A-6��L?~E�����y#�,�?���j�� ���DZ܍nK�bgG@��N�i��W�^����8YC�$~I^�%�l0[������bZ��o:�
���{����0F"��e׭��̫^�z���X���P,��.V�0�Tx������,)�}u���+dd�5��c6k���z�1�(}P��r�PȾ�g��$QG7Ԟ�:�|5.8�rk�:�2jd��t���J6�X�2�e��;TD�Y�i�{�/5�0r!�l�(��b�V1��Vac���� 9W"�c���J�V|�q�5i�:y9�����nf��ag"nLc�ж�6������R^_�""$n9Ƥ�>��Y�̙����ů(r1���wM��h�����^W-q-$5z�b*lE5��M��SCPN�1l��R^F �,s7�}�.�*1�) A4hC��+>�o���l��2��v�������~��v�g��lJ�6�1������I�����n_c�s���sP.�N����I5|T�;�@Zl><ֵ���;�V�P;Ã��8sK��z�r�ة�5t��k�z<Ԁ��@-�͏(�ܾ=/~��7؝���l�ti(��pT��R�Y�ܲ�/�*NH� �����!�3XynXMR��_R���������vu�ӥfAz~�Wt=�|�I�(�Cnȶ�f#�$ Oj���sfu|zR����=�����y*C�k��<Em)��N���3&�:���&d��\@w$�n��PfUd�'%k��ӷN�j"��)>"G]��v�ʓj���X+�����B�_�fT��d�k�^*�=m	�aC�b@�7Y�fH$P5�QkM�/��*�vk;�>�VI�[��[��j>Z}��6�i�;G�m+��)�P)�LY3@�� �����o�s^`M������p� ?��O}EJ)�tߌH���k��q�u�4�N_�Ě>�����'h�;vSN�Y��T/M�&�]/���e�]�|�2��c�4�r��=��?��N����QoNv������(~�X7W̮��a��]���e_
	�%�F��C^���ԭ�$z.��t����E� �T|2�U��lQ�rq1R���J����bɹ[��i+�u<	����g*~y���W���|輟����\̘�|���(�HJ��muC�CP	>j�!�4��g�
�T�'g'�ʣ��E�/�R�������7�+�@���#�>g���;̸5�+�}��&���=�T,\[w�P���z�K��1y�������a�D��ܑ��]��H��r�n84�~�_5�2���s���z�d~E-�v�)�ے�q��bH7ۖ��6G?ָ�N$,�?�@��(w�ّY�WT^H�!�Ջ��]S���傺ϧ����<�l":��0����W�_$��2;/��7�˅�@#~�^2�R��k�|��b2��/��V�B珖vգK�b�z1)�A�
ysx�Ñ���.���s�f,^ؑ����̓R�'9EY��W.���is� ��'�Z�]��s��l.�n-����%���0�CD�(��@�$J�B�H;%�gzh�a� Iܫ���T1���)8w2]�8Z���W�mX�*�NA��>Y�;��o�5yH���7��N����۔�f��`OV��m�w���7ܸ fx�>�޹l �B���[����[�����������ë�6E���(�]�Mh4<Pa�d)�=��������m�ADU���q.wP6ЂRbK+H#ﮆ��,Yf)p<j~n
0�
��M�[��k�����$'Ozx�4�Y���B>])��&��}�#F`t8ś��XV�����N@+���A���ٝ�wJM�\�Ǘ����͠�嗈������t|[S�q��q�%�N��찔��^�g`_��L�o�j��2����9V�H�;2@Y۞%a���0�W��
9�cc4epA�p�J>��o�_N�����Ȃ����fqH�z�)BI]]�lG�Ha;vө���[%�#�d�(��N�^.��}�����-ٺ�T� �%]��L���Q�K��n�0�:��'�������Zu2?����u.�]+��;�aG w�S;��F��.�eM��g��i�J�j�����$�f��f�ȋ9���ey$�������,���oR��G'�_� �+�ѐ6��g��W����D��p�x*��ح�<љ��;��ކ�7r7��ý	�x˷���9W'�� U�����c�3�oW� ���]q������Ź\��#T�iy)�U��ܽ�i�!_p9�Bze�����^32��z�����<+�	i|!�@3O���D
�!�[RIӯ�Z"X�CV��+ 2���2�64� wk�Bn ����⣴��h�wm���f�]{�@'�7��Ç12��Vϒd�*j�t�?s�a�w�S͉�I@���E@�O��d@MexǢi-�n��Li�wͫl�_�AK	f�����8hs�:�Jl�R<��L�XT[qՈ�)cW�IS
d�5 �}���u�z��U���	��{љ���� ������g[�����辡���N��\�n0蓒�:�q~�?aO{4<�o��M����c�_��b𧻓�����;&�E�j�n��K]%j�������Tb����i)����<F���=���5i$f�58�J�Y(6S����Fޕ�v%6ѧ"шK������!����
U���d��j ߂���A�o�K���Iq��<n���8X{AϾ9e��~���ӟ�D��>�'��5�vw�,��Uǅ��(6�G���V{2�s�%���eN xw9�����7�%wdx`sj
��	������e�H�Wv�l�?2�ͦ��"m�/~���W�b��C�o�֖�'�������=�67�ڎ��FD�0�@��߭3�<�=�~$_X�U�k��������"lMt?���-�����y���c�����	B`�]�4�͡�]��}Y��vnf�f1wb��i�/*=3�.��� �8oǜ�~ ��Of��W\K�w#����<�|�Ɍ��yu��4�X�e0^Kd{�C�+�b�uc$�k�0�D���y��u��)C��5���jT8̱��A��s._�k���90�{B �o�:?�9R�~� 3O�*�R�B� ���@rV)�5ŵ�J*�_l-ϯ�Mա�n�4�m��\?��aSR�qw���ͪ�i��AdP��q=�!��]�S���)]Ⰴ�k	�|XD��8���1v\j9���$�vE�������m.:
�h̒��S��M�9����X,�W{rJe��HWo�ҩ��B�8_��O�
p�*P^`�4����o�S��e�E�#���qΠxY�;y���PΠz?�ӜYk񢗟)��4�#�s� h=\�KMi��Ó�k�@��6�e���0*MZ�.�"U|;f�y?��d�"��X��k�X�_�:�,�A�U���JX^�L{�%u�,�jo֟9
'r�RL.���	�pp����0p���Wn@ćQ�c��i�Mk�L"k�rO��d�V |
 �?��ÍR^�؈)p�[R��ti�9�a��� ����O�}��I�KA[n%w��JB�1�&�mU$
�P ���(}�b��iZ
�k�ޘ��VC�R)H��r�{�ƙbfq"�;�|����*l��%c�,k��х�m���/�@��6m�u����=�r���9�(�{�^�z����~��B�5*~�t.@�#���b�H�i���~q���d��}��QY�ׄD-���ԇM�}@���;��ӧ�ŕ�n#���R���任1�	ϖZR���� �)��$���<(s�CLa��+~׀�&M��b�)j�I}�el H�c���^5@DĽ�y�"�%�����*@%����-�l�a@~diD�nZ#��M�j��Ϸ�\�����f�#0n�$P"���|~Vk�F�$�Ś�[P]�;��T�@
+b��uʀ��=X7$R��(R�"ߪ�wJv�H*NR� և�f)"���tt����z���읾Q��sY����<��~a�2�%�LsI)^*����wB�T�<ԯHi��D��o�/$a��#�.�OȄ��6�m~6����)(5T"���<ao#��.F���g�у!ɇ+�9+�#-y�ҶI��2�e��.��BtZ�I�����>��SG�z��y�ܝG$��e�������k��]���10�K� �Áuvs>�G����S)���[F�g���]d���?�A+?d���I�aU/Z(�Z�Q�������B�mX�e�kK�`M��� )j'D'C����Rx�`Y�H�_s��� ���o��P(���L\��I�}���z�N>������j�`&��3���4)Ei/4�	�b�ze�l@�^�(�ƂW���u?��n=:�mKh��tHe��!�5�Jej��tp����ܟd����H�a��奰�(�DO/*�p�6-d�3�1�į��}�)i�KtX$!�n�|� a<�Q�&S���q��zQԳ7�0����$�kx%*��y��}�[�4x�jP2齱ECԅkE%�J�������F���ӎ,�Ӣ�B�<�w�0��YT��f���i����5�roQo.���t�-r��գl����:���y�Y����;a=��$˷�M��#PVR�Kq����å�����-�nm�@x��6݄�b�M�X��>>��������e�}c�FnN���#w���zI�D=-
T3":Xzk�X3R.
��ť��>�q�z��/J$T%$k)ٞ t�?,F|�+��a�I�%���c�v��j-�ʛ��c�1�n%N��Y�0y�ԇ00�����rY#w&���{tk|,�������"m{�� Y��[(@�(C��X���3�M�.���)8��fI9�������G�m=�<kY���-�9gOWQ��&���E�US�g��J'�m$�$y����[�E�D�IO��k	�Z���$�4�kl��;�Yh�;+ʓZ�ܩ�)��v�����`?��D@�bT��Cw��>�#����C.9i��<ӅcP[��kä���_3?۾��?&�)�m:�x����;��8<���-^�#	cw3N&ş׹��!
�4�+�Bl?�2�m,,��,��I���!��)>{�j$�n���-����#Y�B��C�(��K8�����W�����6.sy_8v��>)�W%'�:c�Җ�c_��$g���@	��[�0Tִ:t���*"Mhd����3�\0�9hJ�}�Ǝ_[����L�vU"�0B��\qT�2z���9俎�p���|0��-���~f�n�\��&/�/������ڢ�M��G����{a��2��Im�n�����8��BK�y
F6� �����������-�L3כ�03KB��5��5K�-f��3��~�ߘ�����W�������\��h��?X�o�m�zC������#�2벜0�46��IH��O�����_xIhNpb��y�W�	D����f� B���<ВݔЃ{�Y_�G�eD�d)�)3��hS��:���N��l]����H򱋈c���;g-�f���(��7!��THpB��2��o�a�煾�b��8,�M�fe�H����%�SEO�Ku>��1��r�
,ez���S��2��?�qʹA��V�2�9%����_����q�M3t�6��%�+m<]/����^���0��z^1L��},�Rr���\�p��e❘�Uc"���R拭�d����:�r�����*�.�����ڗ��oD +�kzzj�ѡ��AC��P� c�fRn)2�����q:~}ߋd�Z^&��f�f�].j�ʃyR ����Q��s�1�C_�la����gH�p;��Y�K�{���{���`�	�'(T��x�tC�G����L�r��Րy6wH�vGg��3e�%���ҙp2c*���Ts)v��[���?b_'N������"�NtL�a�G	�PF�0V5���P��Ҁ(w��Ş����82�Z_Z|�r6�_agG�⣍���1V�?���`�����Ҩ�|���t��F�[�zh,˸7#P��ć��;+���GI����L?V
���ٟ�._���D�+KF��I�PR�p��/B�q."v���t8����[��ݮ?�!"��o=NI�����n6I� ��yב��&{�sпL���)=��_�F��wG� �6WШ������G��	n
��&���6(�Q����N��B"���ￇ݌�DwA��<�%s������nrEoEA�ȶ�"��$��kAM{���p6�O�<
O.\��]\����7*�x��G ݺp��!)���Ę���0���T[eU�����8�z1�q*=�!�]s�<Pߢ��T�ה�}������HY�&V�ĿI"����;���e�Ԓ�w�l��9o�����a�������V�@���#؝� {�&�L�+�K���[�q��������XߩI`���
t�Z�n�ۈ���ю�P�r��k�w�}��b�8Eq�����Ϳ��^O��v��dKW��ҏ��6�����۵��
�G����˓�[��b!]�Ӄ�Ҳ_�9|�V`��E�͸��*3�[�9_&(RsoZ�!�0��	���t�ı �����~�B���x�����;u������`Ci
A�V�9G[�[�#�D�h�y���������N%�#�JW�C�шD2!WD+���|�I�]����50�a���z�ݓ<��<��h֓\��{2$��
v5ш�|���Z����=�ĩв���m��Ŭh|��y�y�SS�"�"�Jp���ƁX�Fa�쑱�%�W=�u7��'�N�Z�Ñ�F9��$c��K�� ��ݲ�?yW���}Y�7�1�>�#���;4��Z�Ȉ�3��u�̊O"�K9�e���"A(J��@:�_���t���^|4�6��/�C��/��� ��<���3<��D̜��f�l��F�uy���g�`kyC>�r>q{d���_)�=F�0L�r�E�+��e�H�6�z7C>r��e���,y�����?NMt|ʑ�&�2�"uvO甏4� �p����rU��[�g��;�����qeFl+s�Z 5�=3�7�,S���V3A���L"7Ă�^-���e�H��h�~g>���)��Gǡ��v Qً���2w��fWI>��[�ʦ��)�p�KC��n�ĺCM���EۏDU��x?Va��̇�^Ո0z$�7�H��;F�����jØ�����W�p�Y���a_q�v��Iδ�:Ż�do��zn{>��P��lQ��N79H{��Dm��&�4�p�!���`1o���'A>��$7�[M]d$��`��g
M����� �lX�9~���cMn���?�%1=��j�/>`���G�����>�1�T�e]��4�g$����*�G�V���Q-��
�`�����������3;P�m��8_1lO�|v�t�bs|j�WhL�r���{��
s�X����n�U��?x�sI�/wԭe���)��hi��Qf�Vv*ne��+Q[�8��8���	�\�=Π�#�W,���k���A��+�F�b/n��p 0��|���r�q�P�����9�c�Yo���
�Ph���("ٖr?���nF�*l����q�=xi\�`�(�g6?�-�����Dر�+׃oA��d �ʳ��Lڄ��~|LFenԏА��������@ED���z;X	gYE��Z���V'�*u��ȅ�"?�Tt�-D�����91(�
��қF0�-)!˻*�����Ԕ{Vq��)ݸ�1Ңc��g?h��Q>�TJ���~e7�7� ����"�Zˠ�P�бp5�x�����7.7��}�Xx��`����pcv�#�Eň��P����X�A���yQ2��r6���q�4��u)b{���hs��������9�P���R������v�+� ��9�О�iu��D6U�ߔ�u�{��	i�.r�ɼ�sg(;����;��_�h�Dy�y����2�;�2h�X�hl��q��qW�TG'�6��s�K�p�K?U���w����|���}@Ǔ�Lb�&ZH�V\}&�Q����L�)|��طN�����?�(�r���<G���#I��41O\d)��V"�2B���Q��
������$#:1�/=���*�h�l�m�ۊ�Ḓjp�YG���}��xD*ϑʲ�Ú��@���(r��~M�D��U�Z��w��@ȽL}Դ⍑�<��Y�˹�e� �N��L�����<
��	�9#%����z�r��^Ξ:�P�>3!�W���9�.H�6�,t��78����\�����6�]���b��S]��h�q�=I(`�����3DŇT<H�ZQB��$C"��'�}����*g)��#˕&�w������L��ط�s&qk�s�uw�;���4E��ø�C�������nI|�$c���'��������d}�z�[���j�j�v$�z�U֍	X�=��ȩ���=Yp!������-�uGr�;O�1Oy���W�]bQ��!�bʛ�2��Pʵ׈�a��'Z:�$�w	�ezty�)�}��]6
w*%��+7v�[E�&�Ї^�!��S���֧y<FǞ���cϋ���J�
߿A�|#qe�D�.��~u�N*�kn��{��l�x9_�����/�|�wgxFx5S���`T������HKR�}�M�2���A�Ƃ��)�	�-Ao��_�^Qr,v��l"�r�|-:��RQ���3FC^�Е��Q_;b;{��)�"z�����4��U�GG�9��pP
�[��~��5�bv�y߉p����V.�ET��ؼ8`�Դ�t�02����+S��WXk��u�gh�qT�jv_�->Rw%��^��cDϬf��W��dK����hM�a>7mo�}�q�R_���J��G59�J��|
b������-K~�k/�U1�>��M��yr�i�2��r���xZ��%��� �q|v�����*���h(�ˤ���b@X�_�l&�G*$�/����w�DkOj����2əs�}Tb���62>~,���Q�v��S���	�f3c��8
Y���Q������UY���[�PB	�=��S˵m٭ο������w�V�$�����koS1�������pX�fӭ9�j�Y�@Hf�pL�q��]��)u]�|�Y1���h��=����w�}��H��W/_$��Y�:�	���9�"�@&�>5�Utӱ8w�|V �׬im<\��mժ���_�;h3�:��R�V��P{����ރ@���qJ�}����m�s1�c��t���J�-p�\����śLB����6���������%���&'ui�
���%�Qr@m�
�EwD�)K��&���/��2^U� �?��NGb�qr6�:��}�v�T������Ni��E�m"P-��I����jT�U$��%q��wP!���C�6CYNS�l�3eJ%�-����5_����0�E���eO}?C�����,=8ߜU���܉�seW�L&��OZ����y�&%�UI �|9�.[2�/�œh���h3���g[����9O�����1�Lt�<Ar��DK4uZ���s�(s%���4��� g
s%���h��0l[�s�&(���r�O�ِv¡[������b��03�ۆ(:�������?�#�U��
-Ô8@|
�Ӛe�n�7��P��l7�����a�����5����z������;�q9Pω��[� /ڎ5�N9@+�8��}Y���@k��Pav�e <�x^9�&��/�9L�Ep8�u�:D�qQ�j�E����_�pI^����^%K����P��ȿcSs�\�1��}��sx��h�!'��hYw���(�x�����]eKM���~;��Vtʧ����[�x^a�!� ���^w�C"}v=���y�	1ʦ�eG#8+���T�����������)������R7�/$��x�[wύs)�)1���is��ϹW]s�=!}J՗6;ܜH�bٝ�!�(Zu�莢"ë�5%R�m�6/f�;d���,��cy����e�M�I�= �7�i2����pR��(W�y�(�Vg��� ?Yj��0{ɮ�� 춟���vO! ˢ���M�!�Cs���s�����{�[���y�v��ua)�e��6��z��NZ��{X;0F2Q;�`^.���-S\Qw����AV�A~�̲[H_[���^GP�(�S=cױ��n�Ƈ�Y;����L�"����H���m.tl kf0���-�Ow�]��a|E� �-�-��_�T+�kD8�ؐ�.�Kp��2o��1KK����UYh�X�c+�-e��y�+

���Yg�h?1i�?�<m���W��� ��/)l��c������ϊ�.1q����篞W6�:��D!���%F�t���d<��Fycު]�w�[ۻE~�K��
��?��׭��Wg�$�Crn��Hx���H��bAmUH�L�X�%���_�2�<>z�',N3K=h7 ���T4���4�7���z��5[Ji��$G��NC�'����h�3ȵ�q����.�U N�Yb�]40�$�okGE&�����i�����t|,ǖvL)୵�5^�~�B^�%�թ�|���x�8�Tً��0\���������Ք�B�'�H�1>s�juA����N^��TG����W�����h��a�������F�r����O@*�	Aa���E�m�qv���#�Y� Az@7˔ׇ�������A��UO9@����].�Lu|+r����Oj�h��yT�j��sM�g��*3�K�<��s�k��}	EZ��½|{���y��T酧bЫ�L���:e��������mԤs_CB)Ɔ���v󇆗Î�'�L._.�Z��師Y����y⼥�tB���-�^?V&:uB��U�/1��lE��6�Y��=;�z#hfxba����Ԡn}�2 fu�Z��Υ��:�� ��x+V�r����3����M���[)Օ�\�˷�1Zs���v�l����l��*�s����#*0Gd�o.ZSA��;@��E�X�mڅ:M�%�-��LXb	T"?��]C�gQ*�+���u��hf�~4�힜7��ϻe3`�S�@�� ?�ARd�WҏgYo�h���8�k�ʏ㫎�����+�b♡
�EG��6 ↂ'l� w�@�9��7���z9�gb��Ds5��#�DU�eYYi��-�~ѻ�z0��Uu��_(4, �n٫B��Ǖ�5�m���E2�����q����Ɓ���}��&\��D��a�#b>ioG��F�{&�
Z�ci0�P��O�/� ��75���L���Q�܊a@���,h�zc3�!߄h7�E����5�%��L��ù�0����Ҩ��ہ� �#����1�9.����Cyo������2A�Lr���� �%6?v��M��/�MǷz�eşu�|q�0~f�JPZaVش��< �('��ֵD(5/���sK?�|�=��J/�t�1�xD&z,�H��&��2�P�������ɧ�6�$�b��o���ec?�� T1�#���e�%nU���:���o��X�Gb����2�,�ͅ�[�x?�$i#�I��']%�!�O�w�����0�[_9���b4l^KԂ�+��x������i��i���Ȣn�&gDz|�@}<� �e��p�$N�y���LȌ�pa�]����v���2`
���x���l��k��a���m_xN*�/k]L��%{	�f�t���#z΋tE�N�y������tE�!8�Y�,$�z�ф}sC��W���V�_EN).P���zA�J?N`�AtUٸ!\)�ߐ��uD��?7��Ӕ�z�6�����2+�x1���p�<�)M���O�}+�!�ډ���a.Bu��뿋���T��f։�%��"�*0p�䄇���)ɟ�E)E�������]q��ܹ5,Ɖ�h�b��8�7���5�8#Y�{~ۧ�hX|���q�S�����y��hO�l�EI��x�؞)W�a�_��y��]��)ğ��4��>��5�om'�Xh%p6��'��#RWu+��}o_b�1�D7�l͢(+�d�|�S5��B9б��r0�j�V�I��R�?1m�N�э��l���˟߰����9���f:�O�l2KN����M�@M�j^Ӯ/��xќ� �Q�r�_����O��FbTʵ��A�$�Z/4Ȱ~��!j��Iw�)�X(ES5֚5@�P�d�OHAx���h�
??�H�51�$XQ�$F��W�D�~U��Չ-w���Qu ΃���۵Qٌ�4W�5hy#�Ĕj��'���C.{���(�]����pmze�DӞz�χ�����j�=��e<���A��%�ǧ=:ڍ�1n��1C;��
��i�)mw_���wuOr݄��Q�(%d����+9&Z$0��M��<����(�̯���l����Bղ���͉�`)M~���H�ӂL����v�s�O�PD�Э�o��c!^^�lo
�r;���'O���t�f�A� ���K\�.
*���(�o�hv'H�樔L
>���S�t��V���4��(W��+fx����'��)�)�o��8L��t}��&����T1�p������,�hD��|�l�Ϟj���G'
[r��S`i( �h� ��M5��_��+�[���G�u�<4���>#��7R���D��}`�[ޒ]��'qz�Z��9y�_	*�M��Ό�K�~�g	М�If�$*;���	F��p�#Mj��:v� @���i"b��%  b��8����EOY6e�@O�H��]C|:�P����,����v;���|G�M�E��d=ؔ�T:6����%u���M,�e�IN��r����ȓz������]�xz��,�?n�l�Y���ox#��7�a����L���1�G���r$��lɀ��׈�SS.(.�-�kp���`�P<2��B��pؿ�;bib�xW�C����(qt�{����� ��A/P�_~�Wr�jV�v_g$�u�xH�r�i������=s��*��+\*x����m�$�%��4�~����hb�.C=H����9�Qbwi>"m���J������)��Ď?��0��`��`����V(���^�����o��2C��eF��ꌧګ�a�u�A���}�_��&O�G]�} '�U��Kl쀣�7B�t#P�4�'�%��۹)�<b��RWt�8�-��ׇ�P�Ԟq`��ǖp:����V�31Y��_/���F���9�+�����1�s����*B�/H�y�\���NdY��V��6�aqoֽ�Mn'�p-I����a\o=�C�����f,�3�������{$���z���6"f��\\-\kM�,���Ŵ�1UV�?GFd��ͩ�3�Vs���J�BJ�d<�u��R��4�p�����i&���ɨ�3�.�a�;�x��2l�����?y�����n��c���8k��+�@+�O������[����~�����&�-�!��ɺ���Y��ƛ�� =��N��\�\�4���i���i�q���ݯ�	�U ��S��%����<�2s�K�r"�e��X
�CN�L�o����C���#���^��k�Z��AfK�$_������R�_{]-�0ws��#��i4^�/#�Դ3�(���'���i�xr����O�)���*]@�b�vh0�����M>�+\L�b|��������.�"�v����*j�Y`��<	(���Z�8���~]�����UP��Q}N��]GƑ��e������	����g���f�L����N�eYxd;��$*K��a.�E���Ai�� 6Rd���3��te�ģ��X=�=���:]�Nv`���
P��Z��QMD�x:�#tL�������N�f!Y�,ĸ�:���%q�[I�Ɯs`��<��J���JE��$�x,VnUN�����J4�~31��D-'�"<cH�@��B����^Ns:V���T(���JMA�L�3K�aL��|�f��E&g\'9��D��v_9�q��5K���#胨\��� S�&�6T��n��Xy�/0�"I9VHe3a�B��� ̪�xɒ��i�6�|@�Y9���c�*��xG4�\8r���$C��gBB�z_���dŀ��nZg�/>���顁,�x��ݫm5��%���(�"�F�/޲㯮��(s���_k�'K!�N��_��I���	���с�P������!B����l_y��j���z6�3�:\01�����~K.�Vc��XE���If4�g�.�Auvy.�YK3Ͽ;�W�\���>��|���\fF��,Lz&�$�F�|�3 !���Ѯ�O;�F>4`-sKw�p�K��Xpt$�-�?�6�y��a�fc�oUq찰��لI,8e�G�z����WP�( ���d0_C/�������*y���[<-�x_*�.�L
��z��r(�$��>�k�,��#9�w-��v-�p���NYݘ�#�6FV<������2K��>_~��s�GQ��Z�.1H���u�*.����Wu�0f���%	�WW:�It�[�g�J?��8���>6 ��컫+K�!��Ӡ������b���ِ7������(��j�X���>��m���BB��I�L
�!��!9Мy��J�%�iQC��ʝ��BsH࿰�Q��_�0x�qqHˋa_r���'r��[�������A����2��'VѨ����Q��'��`Z$h�t�y+�����,Cz�x��ϻS녤�LP:Z(�Y'/����߀�燎�p0e�P��h�3��>��o�"�ղ��3�2�5� �BQ�4K�����!:�E�t�@R!L�>hyqߔ���ʧ34���V����;]N+ �:��CI^�(qo����9��g1���C�JX[G��'��u����(G�L��r�H��w7�y�
�QD�S'�&!t���D��
lk��n�(�8�y���<�`R��>��9�n���]s�>������gb�*�s7��R<�+n,�_���D9"u��1��9"����f9 j(8&�ݵ���Tq�\��;�����`�&��J�JX<���8�\��_�>c��3k��y�h����ք��&hz�~�Ŗ�&w04�7$Ha�>vY$�
�g�#X$�p��O�觶bH��������)�b�-6��6�n9c/��0���d��������.#�H��	s����M�uK5s�B)le��[;D2�kY�r�Sg܂1��@�X"��eiL]a^<}e�W���1�L�XR��4zM/<��]YĽ���_�m�虁��ʟH=m�b�?�%�X�0U@^�#Il���? -��-� ��jV���&����{,�CAƐs��v�JHt�0#�N��0������g��.������G��T�N�P�lq�.?_��f���io��4t���"N��?g�Yd�b߮�zu3�R���2��1b��H�)Zc�t�C��܉�L���NT�5��x2+�؆:����?�]�� R����Y?'�cd� q��[�<�}`P4��A�� z$!�|��=P�3���ri�z��̃�D%](����o�tx�ey�ˠ�F-�#�������&Ф����
&����'�| ��Iś_���Nv�3�����0��ڥ���+h��~[i��� ?�WY?�O��cz��-yc�-.<�.�Dm(��X`��*��Nu������H���N�4m)����[�P��3FFAH�������L��1˄����	�b7GW"���9�*/��� �w ���|i�x��h�V<�~���8��b�֍戰:��BLr�b���b<�G��3/֬"�wo���E��^m��o��CT�������o�_"��\��ן�C�*=��x��jr�Z�<I��śH��d�n��y��j�A	�}��D*d�Q
8�]N�Ƕ�J��׳�&��}�STx 8Qs�g�����N��7�[	G�R���j.��gA��k�����â�n��Mzۼf�����0� �Vv��SL����`��Ѓ�]9}�+���mYn�X�(m�B�z�ܽ�QrӀ0��/F�e��X��$���LJ���%ݢ
�5��*��G3�Ѻa�D�O����l�`.�CƸ�I^�d�s�����������F�ZT�$SmA�q��3��-5QR�NI7��[n�VЅ<l�W(��G�L��)���Д4��֟��,�>��:�lގ�#�pq�jM@ �XJ�����7�'�A�	O�}ZQ��K�2*��(v�a��_O�&��u:�O��GZZ�oNVί����IuXZM߆-`��4u�b��S+94Y�ul�jL낚���n�2��7��-��N��`�4j�j�n`G������S �{���qZ���p3�(x|#����陡�L�zt��{��ѪgW�q��.���Te>#��B�nՑ���|/�H8�)<����.�cROk�zl|EEN,[�y�wF�Ԟ�A zق
_�m�fƶeo���τ\O�/t_�|6��W����e����Kɞ+]��!��~��8 ��	}�Q�-�YI[S�R�Qr4]*w�b����W1vm=��1 l%P����3��:RT�����g`,�>�R��a�b��gfh��]. r/F;?����<����e04>S�#���J�DZc@Vִ�[mD�շ�:��a7�����W5������O��uY>����t�_K�^�ߔ]��$�?v��4�M�o�&{����#�>:�c� ;���b��'[�מ������ͻl$�t*	���������W
����R�M�U�=��
��*d%J�2�g��N%���x��h�&1q&탷�P�P�L��j��,�]l�J�L�B5�_�<VC��'��|eף�V��b8&MQ�~=�</���G�P�ð�m��t�󑞎�
��4�L�_�6��{���{�5ST/��[�^6���V~��v�W1�S?�xD�YҸ���ݶ{ղ���T.�_5���XѬ]��Yr�������`p}9��p��2��{V���M8��i�n~|UD̑gХr�O��pJ�CQ����铮��F-ч��ߏ2}@3FbS�yf��k�2#�u^�NH\����ߔ���C�w�/|m*���4׃������M,�A�LDV�A��}��|)sy�:��]M̟����`=��wO��T���)�����X�濪/mU��T���!��H����+lr�Z%�@���q���gq�`��ӵ�r��+и��g����@;2�
:-(����=6���)nr��*A��B{�l���[>~�N����4c�tp"Ҭ��?~���)w񇤌yZ��)n����T8��m����m��i|l3��&e�-�%hlpƆ�w���n��Zہ�2���gMV���� OH�˦���= q��"|g?z�5����/�dZ��K ��{3-@��Px�}��'S���vOɠ�ݴ�쓟��zB�N���(w
��-�D���;�#��������.�l�m�FXwH�C{�H}k��}�/>��	h���S��INl����[�#x�B1/<R�{�f�V��q�ँ�����Y�C��Wp�/SKg����\����oy3�<��t�HۥjQ ����&��
	h��P���N#�T��yN��h5��@��ے�����v8��j�l7YdTiڮ�s���-�������m��Xc��~��6ޠ]4��N���m\��W�⇩���i =|�O?����4�����;�[!�g�4���m�V�V�0Jh�qt�[�W�L�{�M�&˪M:�&�3��_��tV��z�V�kNM����Ԗ2.j�w�XĊ<�2a*,�(�\T 4�~2������Ȱ�y��7}���;�f�O��YN���~i���� ���}�p|�/|=�v)�mf:L/	1��(c��r�>��8�ʓMGI��|����	A�jQ�o� 	�x�Mg�\X���Ce�({ˌv(���^Le��1��CV$���%�+�0��6 �[6�t1�t��(sQh4�9�g�,�ޒif�m�w)%���s��3�wt!Ŷ��f�]8Ss,���ȣj0
_��>� �4�&�c���;j�/�:=��O�}E�-v5tV�kyD�[��5.X�)@�u��T���EGd>�u�^�Q��gҧ�Pr���h�χf�5	R}��Y2�c��Xƍ12�h������|s�4��vR�ފ�������R3�@z�UyL�����Ghi�Ҡ�V�=�d��0�;}ؚ�4r�nq�dN�iA
	�B�[��̥�������D����j��Ǜj�}��]��1|h���J��"Ĉ�*l�I���8t�E�b¡�,w��	���GE�(���8�% ��4��=�Q�iy��6�����@�I�
�5CH�.��V}�o�8r=�ST���-�y�X��Sff�c��.���f�!Xn�_��D����C�P�p}T�M�,��7���:{Y�&�e6�Е�g�6�W��83D#d�G�1d��g������"9Y�q�!�g�D��V�^�W!=1��Lx����K1{��>bcA��G�46jd+a�i�� O)��\��o���e�@Ql���7�B}/q�a�N!�dզ�F\����y-@4��=�5`	^��ڀ���m�iBK�@l�ײ�'� h� ���b�3�*t����qXP�o	��o��{�&�Nkf/]���N��Ť� I�HDz�����G�"�HX�A�B(��������B����9=�St|V��\!G�A���{jQ�vl�a�uӶk�Z��������쩚�[������Sq\$.QX4g��E�!�[�6-��TtM8;���`�B]z�`��ٌ��miSاl������" ��5�<�@�F@���?K�TUT�!Q��&{����r����.�'VbΧכ@T�c�7o�j�4��hU{�FοYI� V����8�Ky�nyS1�
�)�u����y�ʤ��~�s���]k�pő�]\�b���H>�o�_|�b��'(]tTJ�j{��.�{Ć;��zTJ�8�أ�g�2v�]_;�=3?ꖝ���;��n�;��_��Q�~_�ʔ{j�g��vm*n�'o6+��BV�E��PڱR�U�j#b���`2ب� Ǔ�����G~ORl�a�<w��1�)�t�ސ���eUޯ#n�s������lN�Ҡo���3k�l娆�J��C%k*.��+qe�^7�f#5A"9Q��6yR�<gO�Wf�$�㜢Y�[AS�)�8�⟇p��A�^²^b�)Y�2�H��	���Q5�x�g�˪V�+�a�-�|�au#ɜ$�1��MC�����TU}�*��r��YoR�D$Ȟ��9�+?ԫb}�k�|�$���05<z~]J���/�vd�Hw&jU)\�]�t�R��n�e	�8v� T6��9jF�#J#o_v��m�"�{QTU�i5��e���IC��Cl�aX4�B�}W�&�v�BWWC�5�Jc���������/�\�t�WD��R�	f�I-9���������#�L�9Ņ<�U^�P?#K'����D��@�,���XF3�Y���cǀ��^0u0������GR�5Ϗ6Pm�Zv���1��5����rEm��~5NA�J�K���8�����*�e��H�od3������H/6rd܄�oB�%�x���_�&������R
/��� �g�&�����Q�6b�@w���v�c�~u�
�(���@ 6�v�7���Z	��?�)�~ʣ�=�U�v�8�23>�Q�U�ܡ��a�F`Z�_d�BȠ#Ɍ�`��f����MyR���� ��H"�A�O�
��6��5�����&�cd^��v��L�[H��d��ʵi
/�|�d�w�kt��lm;�t�M���5�p{0�\��� �N�l*�����SuE�O�۪ЭM�T>Y�arz2Ib܃��8G5�]�2ƿ4�n�V�L�,�җ({��*�h��������K���b�B��0r���Gu���Y��#BI�cc�HX�4!����fF0�R�.QUv�R��_8f�Z#�>q���O���y�ܯ��SЏ�i�/�laB��߇�@V0�[���x~�̣Hk%�3���M0G 6LZl�@ؕ!���qJiZ �$���h3?{�Q��t���;�0j�ۑ^�sF�w�ra�B�z� ���d�3 S��a7}��y�_�}~�.� +�Q���оO�Il`�Ӂdk�y4n�~u�`�պ�v�����9�1�y3ͧBk�����v��;�F)��Ň����%�2��I����o��$��k`H�'�>�_mIE뎝��Pܩw��� �}� u҂+��9��{Ig_!���A��'�'�gW�{�Q��M�k׬\"�ms��[��{�OBy��Z$�C�ç	o��)
�+q@�Z� J5�(�,�I�e�S�c�;�@�c�M=5��>h7�/ˢ�MhO� /�D$X�87z�� ]�� ��Fs���U��R�+�a!;�����_p�F�8�,_�Κ�8f�9�8�A]̔wo�}�(a�e<�`@����n��ō�����i��@��AJ���@�½te��yS~�O_��,Z5	�]��豁X2�ޓe�$?�Y���&�i��;nh�ζ�N<%'CD�U-+��?���f�_Ċ!�N0��ӥ�v������B?a2��_Z,���@��<�8-�JzbY�:9\�$�1͟l�X�6pa6T	�_:�3w��s �ȑ��!	�b��O�IHd�G������ă%�UY>n���n��߽�D�q�R�4����$��k��D�Ǿ��OZ�&zЃ��� �6�W?R�E�G*.�
���L)y��y�oVT�C�wT�Fla���a)�s�]J����!6I?	,�����s͑��`g�$���|���I_�ئ���OM���s�+��.��d���*+�Qqn?NA��q�a)2����Bɼ�;�'@�B�.�/W���s�ʕÅ��B��4EL�5���N`�g�V$9��<�@7RS���O�CH��Z�7�f @�� �<�����@�y��?J�k7��gt����� n�7~�"2�u/��1K����ȡ����{�����a����Yz��](�Ir��Df���*|B��=����u�5gh��٥�l��[�F����Y�ԯt2j�UXV���}�h��[��1�U��A�Jd�ƃ޺)�:�IT#���E�D��v5"ŞD]Q��Ą��h��v[������8y0G.>�w5��2b�(/��#7���B���ƾ���1�v�C���	�n�<���#d6X�H���=g`%��[%� I�?[�������I9�c>���N��`��sa����$���$��$��^�܊�qb&��E6��ԓ�B*X�V!�\� 0kR�KK�O���._�&��_@��iϦ�i9�� �0F�)���5�J����]>q�v􅑁�`�_�J����s�r��ǡ"	�k�N:n���;�d3����
<���1�Rr�j>:�,�K����
i���p��eC�Q�·:xi�j��,3�is3���?��t�}9S���p6�@[n��L|[�����
n-�-[SիH���B�|�H��5.ۆ��J���̒����[�̪4d�C�'��ЀÓ�DD�36]p�U�=�ݨ9	rr�H}�֪�h�e#��q��w�K��]�������3����, 4͋���X��_ph埒�Y��j{u���P���+�Kܣ����콪S�A��tF��K7ߛ�Ѱ}$����=��o�>��X�+�⾔?|͙�.tW�I�>ACʨ+�m+(�{��3�9��>�9�2B�=�5ԩ�%7���FE����c��WR��R.'�<H�Ӈ^}���58�E�DZ�&���/�xm���0��ʠ^��X���l��5�R�܅��f�������M�J��:L�U��2 ���z�����o�!��|x�b� �Km����s�.����+X"�op!x�k�h������|U��I"��6e4��Q	`�䂚����q�v�Xg͜��}w�����f:*���93�gX)%W�:�\�Z�I������p����^c����yѲ�K)^n���������(�݆�b���p%�'�b+��	���<��1�n^v�:�>�	�S��{ �� ^>{����j�+���Y^e��72���G���Pugʇ`��y�&Q.��'� �-�ĺ����l���>/��ee"�E����%n;9�[]�'���kcIv4���(xcB��ԋ�n���Qʵ�'���O�b}��ޑ���Q"^[�HE�'���)�c'q��v.О��!�^�UQ2v��;:l?�%J�5h\�J[��Q��Tk-�OĶ��z F'�/�o�}�1z���^P��GL�L�J�jؾ�2�%y�$hI����O�-�g�9".O`�����>�nP�m�5��f�ܨ�KL�:��w&��������+$���bRT��@�T�Ί5\�C��q�$�,�CU�É���t��M��q7��n�wzYrHYP�5%���v��R
����`����c�i�vf����!�7����SO,��R�/JdQv_����
]��Ai��)ĵ��Dy�l\tCU��_�׺S��N�L�9�D�����@W�b�;@���Cws�l�t����V*��"WG~HM���&̃�hG���w�X�{��ɺC�Sf��h�"p�Q������
d�J|�0-^wV�Ǜᯞ��A��(�R�2/m��L�)OE�%(����'�|��Js�}�P�~��ц�c���$OK.�[��0+
_��KA+-
oqb�g���gGWQ����*'yy�Lb��:�֭���3#���۽Ř�@H������I)�}�c1�B�g�?|����4�����Q�܉��6E�Ͼ��o����c���A�gO�NQ(r��;��W�7F�����
·X��l�貦�fM�γ	!(T�(
��������%�s�TE	ŔߚxCd9�`?�?zе��X�КU�H��bM��gx�/}���Dx�ƥ�M�g�i�&lF��ope}��wp���F���`��-��;y���b~��Ѝ�Z���$����4l^�0���	�6m[Z��{�[��uB�h�k ;�!�����1�K�h�t)�?���I}�a�4<<�Y��['${�j�S��$��AD|6��O��	��+�o$~���V�"�5��BY�p��y�R���E9WI�賳��Z2����
��'i�fzU��b8�hlu<�	f�M���ً�����mz������)�G�,�VwϠl	��RV0^�)EH4	~����"���W��� �!-�sU;�����h�*8qI����IUbdxZ�jE�^H>���_������g��k��`ᄘ�#���wZm���2㓑��[% \5E��.�ey�7=� ��.|����S=����ڱ����"�r�
+w�h��M�׬��T�+��'��[���m?�!M���;�:ńٽ��	n��'��~��;�e�os��F�K ��v�_lK���S�[���� �����@���;%�EЉ�1�������g!��V�s������@���9�.����k���^�ʏ��T��+�b'i;1��|�L���D�Q���f���/7@�f}���c��/�X!�'�������L����B��<K9?�'�e�Qy�e����g���̞�(���kMɕK���/IT%��4������{�-���K\���p_R]*�T��N�B#:�����L��#O��a��U]9���Ѫ���{*O�����ź¨��e���՟�` ��=��m+y�W�1'�:&�HuO%��\H�s�ӵU����#�V�ka�H�k[1H������R�����&C��Z�u��T"r��v�f��1���s�<qU�Q.J�m���>���4|�(�t�DZAǒ���8�&�k�;W���5"��h��LB�� �[�ʣ߼⠬aQlK$;v�TpP��Ǧ�L���u�cOEp��pN��OL���K������Y�w��� ��Zڇ_pY$L Gw۳w���j:�Ƥ滹z7cO�;7�q�F��i���}��{Ғ��||P�@/N�i��p]l�u�g�-�z����K�|��q�:��?)�ZO��x$�KqM�o�����nsq�V�}Vf������Plaz��X`�	n�8�9�I@ˇ�7��F(?�=�E ~���U��A�a`"h���=����ʓc�D��D�A�.{�F<�-���s��^��*�I���^�9����M���h9wذ�W��E��<Z�%�F�fc�>т���D�^wΫ��	�#�P��E��Tp� ��ջ5�!�'���Q:�>��ON7��q��iTD���WX�V4oC�D��1��*C� g�K?�b3����%z�Z�P�و��#�9q�_�7*8�c�<��fp�/ْdmO>����/� ��:w��NQ�QK9�,�T���J,���m��j���z�;�.�1��?���*��YL���j2�䥠�'#���;X��k��x����c�{��[e�i���%�6n_��ij,ޗ;̆i% �����]�(��L�������ᨮ͎o�����￷s�C��(�:��,/��x����/�/�I2Jv��@M�7L:�y�2����k(͆}y�6��
<�詽�C�2od����rV2�IҶz�	KZY�J$�n��>F�N[�Ͼ�q�;�f4�(�!,%N�c�|�F�ƶ��p�兄siHg���iˈ�8J�F�I���;��c�bAt᪓���J��
�ZY���_��Ğn9���Y�F���,������Ka	���5����2 �4�lo�+S����n?�'�8�1�G,���gC�ߋP�׵������ �B���^�`���k���Ǯ���ɿ��ڪ��:�Q�x�`�1���gp^�L�|K���5V����~O4������ׯ�n/C}u���J��O<�#��%�N����QL!�d���u�{	;v��\>s� U������2�TѫTA�]�L>�@�ܿ6n��r����oC�� �jG%_4�����P�TQ���C��5�	�?hF�뒙!���a"oC��_R��7]Yp��U��4.�bK���+�is� *}NVXY=[ȝ��=�oz�]R� l�	�Z�d��;1ߓ}K��,�>{g�i�wʱ���0&f3�^�x�����=+���f5?87�<�6����ڍ��k�l�)��5����֡��=�r⚤��8�� ��AF,�KZf���U\Ƿ�#�Y�oA�8�'����/Y� ��	$�"ʯ�� �����1V� �P}o�!#��x�gC�@S�w�U-'�X��`1wh�_��I){kj_"�'�|�o�|3.K��S�\��y���7��p�ɏ޸��6�{u��ym %�<G���RN5T�p�h��.j��p}��cj*�����tՆ���R�S������4�ϖ��rӣ�3R���'O�M���2y�?G��ү�CO��"��0ȔTN��Of����S���t�Gh�ك2G,����L�����֖'�Q'����{t�<^dDְ�*��5�|�S6W����㪍����!܈-9Ι�p���R����$����H� u&q�~ ��Z���PS 6��O&�|9�VU��k�pf��]��9��av���.�2��Ӣm���ې]F�o�s��is��G^�z��/������j��[E�P�R$t���� �%��~�h:��[J�ӄg�.�~,�1�x�����@��_II^�W·���{�X_��W�|�ޕ�P,U��{���-�ڋ�J1����#	����i�*A�lE�hV]ʖ�+23�N�)ѝ�݈��\���$����&����~Lx��& &`��}U*?<�����y�t\���z�۩�a?�E%�⨗<����^�c}�q%5ķ���_�c�6�P��P�y�ʌW����+����q�@^�"��F�����n�U|r�[��%��n�	���+��iC��iC4/���_: ���e�d�:�~:ܨ&�y�`5�$�q���< 6�`q����1�ri1�\ހ��h`mA��Ȗ*���'�ӛ���?�m����J��=_�L�����nkүP�,�1��w.�'`͟�Fw�$�� K���2�5��,M����!��4��:���thI��֯I A��Tf)����E�;�����i�	���:����}T����tc�Xx��JL�𧻫s���Or��
���6;��Tx�1#iG�QilJz+���N�5f�X���.�{����\"����z�-PF>O�e�a@���,[�.�#y&0����vW�N��Mb�TYكX�O~fӬ��/J�����D!����^�U�(��8]=�x���m:�sI����YhF�����#$���t[�=Y*d{��x�Z���,u�Zl~B��j+쁇��Ui�L�N�h��f���Ӥh����!��~�k.�+66��a8����X ����&��^�U�>��6=d�D緦�;���|�08��kX�e�	CQ�:�V��4�	��fz�-�p�X�#>����ݣ[��},�������D3��T�� �(i�y�-�OC��0��>���{کj��v<�=���i%d*�I!��ts˔U��-��Z�pou�����`��;Q8�R��u�3\iAE�ea��W�x�3}�ǖ�+�Zԅ�|����H��	+iR�^vLbE��	O�߮Ӻ�xs���$��%�*��Ӂ`~,>4G��ڜ�-�J��[jM��)���j�I��s!jۖ��L�����!(�
�:A|l_o%ÍRy�M�8����D�#R�<L>H����K�*B�:YJ��DҟaH����������l�23M�]M*��U8����������8Oa}��c�騐r���%.>�INjw�@}naZJ�����Y��{����L�	���֋�K�S�,��9�,�I��`��֖3�� Bę0�6l}z���I)~��`�J�h0(�����$��c%A7H�><��hmdv�;�k�JoƯ7Šz��hp�/���ȷة��N��D=a����?������
e��@
��f�Nh�M��7.vu(��G�S��[]�E�%�W��Ƀ����$��˾��A���ߍE3l���e˝��zi҂p�u��o,|�����r�)x3y�Q�l����D��H,�N]��5�Fvˣ�#�c
�.�D~�z<�5X�@�^�=-��k�X%�AT-���5�lu��_��Q,��l���'�7�:;��g4���U�7�R^3�KSLcI�x��9�^G�����������^!>���ōc��.˒Z��hiH�m�*V��w 8>|N���p�ȲH�#��ܑx|�?��2=df�ҵ�JEh����:�A�t`@l�66�l�7R�%�;8�7H���M�t�7>�<�6�ʍ'�䖥կ��e�4a��L{��;�j_�m��A�|����A�U����cI��o��6�;Մrd��e��!�$�_��������	����z�x����nS�WsUon��n@����
X�ri�0��8�\�6/��  +�`%ï)�#$�-�.�.� ����WܷI}7I��W����C]$u ���R�i�^Q!if)�=�\�hM�?�����2�i_��/-���woU�dp�
���,-��J����ޞ�B�����v�����;�Ĝ·˨Ǿ8k�LR �G6� �*m1��Y�vcEcQ�������QC��no�3>�����:�ͽd�3�`y4�����F���O�x���a	��!'���~5g����۠Ռ���2歷����zW�Ddx֢l�1�P^�0c�U*��K�K*6�/@SgD��ڜk��t��������O�h�Z<V�T��"T�i�_l��f�5(���]�F�o��v\�w���,μ���䲙���zfH- �Ǐ��e��љ���U���g���
)=�)L����00@�}J)�:?��Jf$0e¿�ߎv>�׌��p�$|}t�� ����F[bu������g�%{�z�Ÿ��R��;q^��ןD2���#��r`�8��-t�e��o�\��y:�vEC�9�C��{I=S�|�Ъ�0+לtÝL#��Bp�L�88su����ɽ˘�}�V�+\�〆E���9w5�3Q�z��S���Ps��ג#袼���	B[����QU)�G-M�¿lP`r�������ez����/|%��!)�<�0�q�[�������(�DJ�)qj�;�u���N(Q����%��*�����e�{u �ƕ�v���,�yo�찧'��J^�ސ!A�fk�H�>4�|�N���
<��2U�؈Q��{�q��y�Vȅw��D�����%Y� MP��ηkQ5��eL?�7$Ǩ�}^*�������W��~�Ի��㬀-������������y�d�|!�%Ԏ��BDxaG�F��f
2��˖��^�W��:��RmMS԰�{��m4;�������ˡ��~��Ҫ���B��R�M�g,�, oD���UR���D�9�)L,Ȍ���8��Z��I*�<���J�O��)Pn�ubq`�#qEӚ�tPɂ5�,�zdu�]�y��\B�l�F)R�u5�H�]��eMt�V�r��Hh�,a�b�gHX�^�D��ZafWPUP
.G�A��3��wE�KO�Q�����1�ۉh����.�Y�N$QzqML���p��˟eb��WUAd�2����҅E��짡OSX�Э�Gt����co��4Q2&�P
\���m��-?;R��~�V�7!�I81_���W��HVˊ��I��Tz�D����1�l)��3�x�L��ݯ��v]pR*�CS�͖c��զ僁�@��&m^��'TJ�e�NˀPNshmm��Y�c����tv���ک��o�jE��_�����F�-�1���]P����Ehڋ9�vB���[kJ;� �(��]�������Ս~m��l�<h��h�h��֏+�~{��ǵN�:X��G�'�`㭉+�!�U�2��eY>2��;�4`�L�P��fs3emEV9��O����q�D4�tH����|
�.�*���wh��{-��j��Y}|�1|��{?Z��ik̸��߈���x\,.�E��]�1z.VXYVrH�s
�`U���kM9a���&�aRB�ްǈ'�U�0�텭�v��dgGj0�P۵��#㢈��=��z��$�FC \���ڊ�lx�@g�1����W�����[�1]�����䆟�K�U��/�FQM���F}�g��mΞ��G?O��}�+��y�
�Z�MR�f>�2k�n������k�yy�@fsH4�����@��$�~��
@k� ��\
�@l�&>�$�N�7'�"��ݑg�:���Ѻ
Ah�\PY��+���#�Cs�7��--��g��ؘ͔�9�i聃�ҍ���Fjb�� ۥZ����b�/2�6
0��5��l
2�)
�/\�x$�n=��m��;z҉y"��~� ����I���� U��~c�]|%�^��q?b���u����=�Lf��v�&�`P���A����䄖@���5�U� /5����+�Ш�M���j���>�1��K�19�k�dԀ`z��Ml���A�t��zs���'��:�[S�����-MJL��\K�3o��@����6\�\��a�Za�4�=���'H<�([<y�$;m+�k,d�r�LӾ������C8h����ts��x%��t,
'�K�j"q�:验��D�Tu����o*p�g:AO��&v���w�Ώ��]���ڗ4��� G�Gn��.9��M�G	��a��Q&!�n��X��|�u��d��Q���"�S�1|�:�+���v��x�-��"��о*�0�����"�h�F;f�{�h�Yh2n	��%�0�x����聾jRWr�2��f��lX./��B��h}31�Fb��٨�A�)�҉?��Yɞ�;���p������;Ϻ�����6��Y]��<F�4��:�հ9c�&P�Ban��9���u��"B�с�T����/[�<��}�Zu�j��ݛ�����ԙ���z�E��wv�J�\V�O�d���wO>���ש&�`e�+aQ1�"�c8�dN��ס�ȐtMӺ���\�ѳ��ǚ�7�y���@����"�b1v��8M�;��g���$]e�C`����z��A���+�KR*^v2�w�O�(u���Y_�۾щ��=AG`���/ě��ʩ-�?/1A _�p����	D���"�G�(^j��<��Ɣ��0�U�
:��J�1
����^k��j�]F�$�si��G��U��A!,�-6��$�Ѵ����VA������mA��ߏ�=�	���A�#�������F�c�(��J�x���'m��������Ļ�.�s�~-ԙM�JL�+|����\ *�kb�t�M���\�5��9�������Z��e��3bn?Im.ٿ������a�M�Eo����> �У�èݟV;C��Ժ{��бl ���Z"F/V���V%�L]?���pHD4�Z1�'s��$��o�.�s�_A�H��/K���794$��|b�~K\Bcs�ӫ"8C���j�r�����In����{����+a=`�Ӗ~p��������n9i�M�]�m[��{�P�(�fJ��O�n
,ϻb��^�:4<0u���rߛ㕑�8��6��.��>���T��6����Ҏ�!�#]V�b�ѱ�Ym�Qr~@;�ـ4#y;t��fϫ�� �4� ���f�%D��i��wգ0���c_�{���M�9spjpTꑞ�����������(_�O�1jX��C������<;}�"�g�F�u�&[�?�jwr!��LS�p�/|-`����~9��������g�C�2�~CEZm�$��˺Y&[p}�-'Wxr�᪓�-\�ht��^$��2ʻ�;�C����ŕ���Q����*�I��:�Z-i[ݬ��Z+B{�(�?=`�GE*��w9Ӽ��~.Ǫč��x�@�	d2�-K�p��(KNϻ?����^��<?��X����?K��C��L� S��웓
b.�T����(>d��Q3ӻ���-�r��|��bx$��g��򈽱^�⨶�����wfg�D3l~Ȕ���а�`�3������5�+ La�a�
I�H��YaI,�R]e
������\b���|i%)�#S�QɇACT9��E��k��m�}���D׌�����R�����ѕ�����>w�7��������^���h~������D0ŋu��{.�����T^�fD�2[�څ�t8'N80���I�M�n�� a!��S-�v��DZs�F�gc��iG�!_�/���T7xV4{���?�����_f=iH�����hg'��y�tp�
�W�L��oz[r[VB+��n�#ogqwތX?Z����&a�a�d���{�I��[X::!a~���zMd��g�ҭ;��dd�^�����7��"t�NnI$�{+�(qDtT2��|�I��IG���0K+�2@?;��*ދe�ȳ�UH0g\0s[N@I	I�)�0+�A��:�$�5�7NZι��ڄMrH\�j�$�i׏�i��Nt�Jn����h���GÔ�}U�x�)�`�c�<�=�T[>`6��@w���i|n�� �#Ѷb�t,��9Z��ۏ����ES�[(.�(��٘�!=0�N�.�0�q����	^�p�`� �Y�}�:�n)V���G�j'�Q.�+������%2ijځu���b�9�a[N����p�V��;Ql�W5��q�H{+!]�}F;���!i�}nd�_o�560���;��e1�*�����`u���^����]L!	�8&%UmM�U9f�0lל�Z<nJ`�?�1�5��?�ڋqtؑ�{o�{�6�4��L���	������:��	���eժ�a���l03$FX�OI����'�fa�e�O~*�����?��#��9���i7�@��A6��s@:TZ��	}��󉠼�;����$m9�n4�j��~y��Ǩ�as.�j&����dr �T�Z��bQpыY�+�ɒdP�4"�3�C͉���b1@y�s[�]a����{0^d���{���Y"s�lM.���D��;���Sr���Ge�$�kJ�/+!=�8��W��akJ�h8.� i>�S���-��V����J�\��6\%T�옛�`�������c�(�`Ȇ�'������le����sg�7�v����a�d4b�Lr51�feՋM8��0<��I�B�XX�k�G���-�e:�g1����}��<�^��P�9�Ӄw��&�S�F<�����館`+�5 �Z��Y�
�!G��0��rV���$�6S�i���$I�s�`��j����_.�)�W�h�/�{<?5yI16<�( ����S�o�_���KX0��� R��U� /�O�&��a�I�7�GV	Փ�i�
l��)1��b )^�������& U-�����1��E�wVȘ����*(p����{֪��:������1�dm��)�(!��ʧ!�3�&����F�I��=J8B�+X��e��b%���B�ʆ� -�:;y-�ET��5f8��@m�>�EK9Z����g�cF���F�˲��·�GZ�<���bkKS�p��>�9clƦ�u �8>�0��O#���o	c��6^�Ʒ'X����D��}Wu��)�i��N����ż\,�g��ս�rL�s���!<�l��DjL�� ��v)���"F���ݠ*��221�X�5�m ��t����IҐ��XDó�P)~c�`�K�U���B��Զ��ָ���"����zg�6�fqFj���Q>�sa���Z���tH����"w��� B���6�b=�Xα��>�-S�5s�9�z�+�C\*Q���"����C�}�7���Q%�,�Gi�������'dO5�>�����VeR�GyS7��������Ԋ��/��.绪w�Wm'�G�F��kLw1�S�?�>�f����ӿ�\��H�/�y���V�ÑS�{��?�d&���ؕ�$�D�E~��%D�2N:����q�π']�~�߬P��������u,?�[�Gi� 5<���]R�Ii �ZT_��9	�P4�e�>���
��dZ�A�*�S ����W��wRb��t�\��]��}�S�xM"8v�m6�J��b��A�۵�y�A8�]��"�z|�����6.~T/8�o�U�u�5[5V�>
�X��c��P8�Zh��C�PxY�Š�����î���&����\U�aX&����T0U�t����mmD�,"�/�*���$M���+_�����ʅ�~��D�ߡ��k���
��D쐩�Џ7�3ۦ*����"߬f��9�?������D���h�<(�(s1QKJǟZݯ�%O���t�[�)��z�A�\u,O^�#+p+M�#�}�d�V�htQtvO_��*W����@�Lǌ�$9'ƅ��tҦG(��$)։�u�q,��\�Lu��}C�ݜp℉[��L��`�敻_��ZjQ[��RsF�SЀ.����C͔|mt����Kz�����v#�m)h�zjzR�lڝL���~��j:�O���z����W���������*5�nZ�u���A��T2W���
,���X"3�`���?	�eN�y�!7$o<�.�	 �i���4��L��.�@���}�cUZȇ�[��lO\ (ݿ�Fi�?Y�Zz��iŝhPe��Oǜ#ʮ-մq���Ά�,mr1��A��H.����oĿă�w�"(�:�-c�r���%����8�H�ܲ5E1*��ZA��l�����d1��O��jۢ���+��ш����J���ج!�G��30f�~K2�X�-y/.�HuFJwX�����c��m�@�쐭����A(�Q+8&i�#�Ж�����E[��F߉5��+E�Ы��äc΅�U%�]ui�b��`~��3aXU�(���>>�@�g6�	�_�+�'��L�eN� ��N�'��$�{��e9Q�ba���D_c���C2�|��T�Ab!}0���e����NK��p��Q���zC/���0���u�l\LS��sc�H��5�Zd����������;�l���5j���jK�נ�=�U�[�� ��3ѮaX�HL%�*��7����)�8���{�Y4��P.�tBi�A�^l�� B�}I��k��T47b��^0ucSH�-⠀-u:�'6V�Z�u�����D��uv�2	�~�Z����ϋ��.��2�s`�u��OvԈ��-���c1
�{��<b�y�W�T�iv��Qh�	�F�����"[;�
��ڢx����a)?�*/�.�-��g.���梞�������b#ҒYi(~���(����e�P�L�	Bc9|޳Lʥ�ͧ4W��|\+��O��j�|B�;�}�K!Oo�\�r@�8ղhB>v���0�ѫ2�\[Xpக	_i�����D�&��E,����/��߳�=s�J:�S�!}~�ߖ�py�)a+�+x��t�	����;�.\1�K�v�AD=vU#ش[4 �'���$t���6��{l=�{_A^s@^�o.�4W��D>�y�}���{5_��08��G;������`Y�3��;��N��G�������<o��7� A5�������JWl����L�H�R]���Nj�T��*���#2885�<��
�z|�P{��>�|�����ϒ����,���4	b`�����щ�^�����)����[��Տ��ϖi�0\E��?/Fq��u�-�]���=�ʩ�o����.�kCO��b�D��Hý(�g�<�����9H�;f�U�ّo�GT�Td^b�BrS�`&���D7b���U�,����|Ks}��������ҳ�'X�e-���]�x�!ǴW�?O��!�={b.*]�@=Ux����q	����,'��!�I���Ȗʿ��̎�[q��,f��.��$���'����쏶8��3�,�ɽ|�uGmEF/��D8a��b��r�|��'U�?�L)F(l��%�BA{��x�s̱���0��tb�W;^�KyRd���)1��W��l��j��+l���>%,8�9�?|��/g)�1e����� a�|1.�LC���#X#O~g_c��{�_�:a��Ί������E7������y2F���r�W���
����<h�N��������dq�[�6}����oYݪ
��:�C0n�W1�,�IFKp~V������q^i��yZ��"�ol ��NxG�2vPg�;p
�3�81 w /j���O�,�2��1:�A4>�W)% �0kr�WP�ݝO�ْN��D�Ӭ����NJYm�9g�%l0Z}��:1��kr(g��o���?5��m�m����Eʂ��䄺p�ѯ�����sfL��,�v�o𷃉L$�&�=+��OR�QE�pډ�:�)�dn�{����p�@�߾rIn�~F� @��X���T�j�B�����,��f6���>ǝ��+hѫ���\��v9��a��|�9��qb����;�L'�_�/�.�	�i����3��.�v�:��L�����l�@=kV����������>ZR��������9!?b�p<���3��t�A���u���F��Eh�C�J2�n�o�J����{�K����g%ܾ/a��=�d��˺4M��'\R=�g������w���p�����-u�D�vD�}������+��m����Er�͓�tWחO��ӯ�v��-p���%��&>�K�x6a��%sV��>&�*}vF�H3��~Ŏ�;k~\u.����n�}�J��'G
��4�� s�dKe3#//��,3��9g�r���*�ۿxR2h��t�g�#Q6Po2v�����}��)$Ș�pGm���_�7o�k���m���V*{�F��fO�缯*>�K���n�=��gW7���O�8�5h���Qb�P��֟������8�����QٽSg�wK2��ȔMz�Q<�G����z���㽓��ʲ�Ě0��r��/�И�"��E��k?#�թ%A�)� �� &rH|�uh��Ǡ��	��e�$-��0�M�0���)�@!;�����Wi6�d�-7���Q@�I䬉Ay����{�^�v3)_����ҁ=n��=ψM��-]��Cp�8*XG����ѠL�궕�"��v�9Q�8b�_: #�ـ��K{,��9Ã����\g�2E�>��N��X63��/Z-�����3;+�������+�\�c��C��W��=M+>�
j��wj�,�,&�Πl�%:{���"�4g�t�2�JKd�=ruu�^�(�h��m&Z�C�;�ksb�}�)x��QL2J��V`K���-����B"]tM���}�rWHv��\¼��˷��;�u=1��nMC��R���f�ӹ�B��?d�s�@[h�����.� O�(d9F��t�*e�H�T��X�T���U��!Um��XS(�cP��?������3o;_e�]a�S����ȼ���K����ll���Q���Q����~���Uq7/�$�ҁ��7j,�����>�7�,RښO���s1�*4�`��SK�b�Һ��.��&�sWn��a�F��*N�Z5��0S �JyL�A�K�_ht���i�C"C��q�a���PC�X	�����pky""�S^|}Hy.��R8L����M֖=��:]t�������qWN���<�5�Yy�q9�.��%r�z���4BN4��5N��K�(o�>��nj�U����OFM\-D��Y�T��h�e����U�t����e����CRV�����.1��<�*q&B˃�Ѣ�M���hu"�=�N�uX�
W�ڗlg��ǟ�Į��x�i�K���֣�+����{w��Ξ��C��%Ԇ�vBT?>Y��Mv�9��/�0�&�"xI��tlU�'��݅�-T�����*.����W>�|R����ӑn��V;ك�%�c;�Q���m�ϻ�4]hp.�������U�Ϗ��O����DP�n��ja�d���-�!�"��M����!�C�_�5�Y��v��Y��H�pRRL�p:g_�S���6D�1���1�&Mn�����a�e�Y4�%�h�=���>ծ�T��e����L���<G�GKyʹAIHC>���N�1BH���x�Kt�^YK�h����q�nULA?F�U<N�}z��?1oL�|P�h]4^~��IY�b|ס��#۽�ݗ����0_�eU���[��j�sg�{�Vh+�'ε6PV'��Ӗp��k�0_ח������e�H�U𓱼�� ^��/��40�6�r�l�.f$�l<e݅���;O>x��Gh!Ӣx �_�N�'���e�]�B����
�س�X*X`�QFFETP5g�����X�U��Sؾj����TP]��)�y�Ǆ���$��ih�޼��索_�n .��³�)$�����Tܔm�7�t���a���S��r�C��Y���������+�:/��Jҷ]����C��;CU�Y '.#1E�~`�;Ŵ�K7���r�y�C�p|��W��'ƗLӰ&�p����V��vJ]cLӌ���H |?�_)�ޔ����:���i2�X����?���z��K����:k�7�[�e� Κp1P_$�(������3�{�L�T����is6鉀$��u[!�:�δk��u �-/�YY��;xIaEOmҩ�Bh�%��F�%�2W(�m�ret�3���+7���j[�*Դ��P��y� �k�G9�3�xr\v��b@�atmT�R�?��×�8S���9�:O��X�Q�Ig�@
k们Y2���n>$�09,�g�2�I��v[Z׫F��h��@��ń��<��x!J�x�C|[���/��b �-b6���wNdE�8�LȮ�2�ġ]�T���3T�qBW¤�X�:W���2�"��.�';���i�F+%��$�����9�����˚���)�珴l�%��I���^��{�~��D2 �=WG�^iLF(҃t��4Mf�|�l�8��K�������!��6���y���A�5u3��Z�+MJ^ w����`��5sĞ`�RĹ������'�@��X���K��c�b5�-�N�Ę�FЈ�����_�4�L���Z�yp0�3<�,3���48�|_�M-������������	����lo@�/�"��7�T�C��P��Zݲډw���jC\yW�_���4o�z��G�i�{��b?㖮�$�q��P�,\<-�#���&��!e�\*U�/QY.!Ʉ�
��u����G��b(u�X�p��q���$Ȗ��O$����G,��"�Z-�����3�]*�yfm~�(d�� a�'��zN��ĥ����O�ے3�GȮ�B �&F��OI͖e�6���U�֚xN����� ���"��t�u"h�2%ו.�݌�� 83�QE�W���]%��A5�!����W:�f
��*j����F�����'/�;8f�֫P��:ɇ,�<	e
s�K���ad�d�Jt��Ƌ�������O>�6Ԧ?��qyp���Qx�=$����E�w	'�T����V,zXtI	O�r��3Ѕ�{EZ�Ob�}X��b����Y��'.6�[��%4�c��(�E�5�kEVƦC��Q�#q�9�>�{<k6�P1���xf���([u��z�,�ڻ��׉�����73������#��5xoF?%��lsBl���,ƆPG�.�sh�h2Ş�"낪�Ψܻ/����$�Wv �;&��#+ہ��t�Ki��6fV�
^��l���$6��Zq?��\�n�𯷝��P�T� ��b噏ט�#a](yk�hHL^���8��4��@�h���jj���c������Ƭ;�=#�
���]G���yO��JM�Ge��#�=�CF�5�^�q��-4��t6-��Դ.^�[P ���P�ޢeި�.���*�V=!�b��h��f��C�e3n�Ǹ'��8�8]��|��i�:~�'�m�'G��O���@˒u|�͌��R�����υ]
��T�Ҝ���'� �lW �9��_�YTl��HKf���?��Q[&[��`�)z\���.�j��K�\pF��a���Q���SF"{Y5FE�,�ؚw�%/�sO��Ŀ�I�K��{�s�p\V2��1�����R�dOi�X���|9�3V)}D�-O�7K
k�OU�M�g|8&�2�7]��d%��+�j������*�_ޖ�&��Q.��:��Z!g%S>Rd�w
yL�1��d(���Px�(s�~�0�Xڲ�5�pd����lFt8p�Υ+���������-_�_���@v��2F"3�����`������ʽ����@C9�B,1�sO�1�Ҋ���W�]JZ��o��y}h��� ����K���(�
h9�ȩ���A�bGPu!�#Z	H�k�\�"4��yWR�m�1���7W[�hïsA'�ZR��v�
�[�����]̔c�Ҷ�\H�}����J/GH�l꒨��6TIHU�_}��6��OYYW/{_����{�ᡜ�<nte*�Q��F���a]rI۟Rq+�A`���Ff0��y<��F5���2a�D�(��t+�����In�`E*�������zכ�`�ҩ|��z�]d���j�9���O*��)�Tq��$�������܏6mŋy�4��}(��8b�.��̧P��`�=���i��N�mP�O�&Gq�ˉ�eVk	\�@lK���`�LqO8Tzx�0���2�S�?�s�����s�r��YH�:[iw|�-��Q��w��6�.K���!����	|�O���KnD��W�8B^WY��h�+�}�TS���B�$�Px�����VI�̸V�Qߡ��(�HN/��	Q�)�F9
q�
/ri�eWA���k��
��]��
]�&��ޅ�A|X��k�\߶DC@��XҸV�� ̉�m'���? Lg��x�7�oJO�A
�������K���Ȃ%6E�j�+B%��zu�T�Sv���f|j����C�!~�>?�����'d�/���pf��-�%�G��+�p!m�>��$Q��O`��k�H`�K+�̷d��Co^�~�O�3$gh����B^*�I$�3"V�-�z��G0{�&�s;��i3��'Y��}����>��<�izɝX|G�X���-:M&�ޭx~�������<�#�+�Zr���Ԏӌ�G��a3XKX�-�cJS����p��?�"���m�Z�s�޽�'��zo�o��"�y����L�4�d���KHc4��j���t���'�(''�aN����Χd;Rz�a ��d���3_���H wWL�A8�z�"m752) p?��*�~�뙮��'���*-��-�5tV�G��}ث3�	?��Q[ƅـq���K���~b��':�HM��ũ�܅7��V�E7F�3h�bYpW�J]F�|�Y�d\,�{w^�ߘ/�+�����JQt����[T��rh3\dD�} ��(�%j�Q��A S�1J+�,���| �8a��N�99m�o�f�S�J�{��vig������Kքy���Y�(��m�F+��H���5It?^�ve�o�Y�Ǣ�r�<f:Ш�SĬ2��S��{Bx,��W���k�sC&��+�L��)J����{y�����F��e�]��^.0fn�4=��F��6E`S�/%���G/�$�o�t����i1�M��ۧ���L�
�f�S�g0���D��w����8�FF4�:�U$��+>�|
�ב�5C�<�T+8�7Н��!G=+Ō'j��hD����E�9N��A���^蘽��M���*Y���ݚ^�~��qL�G�*Tޑz��!C���j�v�����'^T��"���\cʄ���Ҽ�:�Z1�֢<P�]�K�l3�DQ�j"�W�iQ�ȇ{���Z��$�7W+4]�x+��,�K˧��Ԣ�`E��W��>�&P��+ͯ.샞�}����0��j6�)\w{N#�TF})�����/Q|L��\��+�͠���S%�(0�8��։��@pFK������g8�!&�/������zxtp@\*r�B�4ir@$�0�7�,�oBx��_���>0��@�7���L���^�+�95���	/�-=��Q�IP���Ȫ�d����T$�TNs*ǖ8�349��n���M�n0ˀ�E#z{`&����i�̿��΅M,��7��7,s����J�&-�J<+���u��SD��	�q��Sz�W�E�=��L� 8j����fѡv^kj<��Ň��yj^�ψ��C�q��/}��|�cJ�O?�(�CG� �m�ΔPeW��6^��C�h�ϱH�m� B$�{g�w9�M݀��x~7
�C��b`q�Ϯ�B��U��STk�	$�õ�W�+6N�V�?9s�Ǚ�D�i7ۮy�Ӈ�kp�����0��bȠ������ 8TK
��	��A�_�z��jL�$g��V���*���hP�[=��7���� ���pܛ��5%K��������8	5_2j�," =��
�[=�2�������S��l$��Ft�y;h5Mwn,{
��)���%�1g� "���7�.��o=���ގt��[��_9�k.i�A�L\�3�u<2�� ��"��6��	��~�hd~��Y��~D$e�X\�XYD_��Z�a��?b�Tm��re�h���1	!L"�b��/S��5�-�����f��F�=g:8��ⲱ�G��Ed��q���_� 7�s�ƛ� ]��7�������*�P����?#��i�D��(&�������
�	x��p8�V���%+ѝĔ��I��f
��ps�����Sew���ɼv�b��8-�/��"O_K��y{�U����&���~_L)��x���v@�W�"�o��R1�����9q2^�� Du�v����0%{�.�k�ɐ�J������B�ݬ|�#M�S����~3�-(�ｚ%��o���`�E�Z���Y�_Mi0u��@����VF9gg�7�CY;��c�fnO�n��Vб�l0GkA��VݭP*�/k�a�̿����㗚q�<�է�R��������DڞHm�s��cC���`��ƾ�b��*i������S�j��������1�k7��]~�21����>	Q�;�܊?��ؠ���+�2 #:��sR�!g�}�L9;(ڝ�cLp���,3��d�x���%E/Y��=�8mm狔{���<D�S8�j�;^"���j뛚�t��`_�)s�>Fn?���>K�s�\�t���O�p���Suo��<��хμD�����L����܊�x)QJV:w�Ԫ\<�q�QG��I҈�Ȅ��VG?qjǺ�V+�:��2S�҉��r�cY�pH��zTν� ����`�A;�q��2s��d�� ~6��]����"��#v����[@�Ig�N��]�p�_7G�����/�����"!<�t�6���Uy(Id�[i��iY1��VnK0v�6p>�76�r��W����4����<a��̛���Ǳ�\u]�D��CJ�������C0NeKDk�>R����ٶ4m�C�y�L�[�[L|�YB)0\$��'Jy��������"8l��\�Zo��-3��Z�|���D^��������k��f�k���8��j_T�D[)3J���Re����
�gv�U��Q.7��<L��?F�'6���0�vt��T�(1=:$�|ٰ�B�v��.�T!�+���`<�)˰\d�C��Y\�W���6���	�!��~��w�-50�dm�ָN	��Ib��gW�b-��E{�\t�b�����xVlK�<{�����B���tB����a:8�0d��
��&]E���`'��K�,�D���.��;6�kWI��*i��!Q��l�Ķ�#���v�*U�E�8�^1�-�o{�N)���3����Hl!#�#��	 �o�gk{��|�fm3
�$k����,˗װ��������º��#S��޴�kv���o�ɋA����_��P�,�Ǔ�@�(�Of�l̊^����x��$�u{W'�NG��@l7��	�k�郝{U���o%�������#�g~{�n��7^�oF�2����yv�[7�V�B=h���ȘX�fx��2x_�9R9)5�Y(����d��ܠ���u��-�^��X�Ye��x��c\��R���~^~,q
�R8��?�2z��YZ�R����T-��bt����c0�.ޣ1��N۸$O.�0�VS0�m�
X�pJZ�%��j���<���k�����Q��4���;6�!PBز��4l��l[�f���+��Z�q��1*���p$��d�u�{Z..)']�{�g�kv��a��2%p��-��o��ܸ-ߒ�0��DC�%{���:Q��Q�����5������`�^F_�B���M��� <�`A�A�s�:�.@z��BӸ+m�>f5��������q��9'̾�_�g]��� v�o~��R�����q��[e?�Vr�s�hnC��Vܽ�O!�;�|����C���e���C9͋<�3<�b�P۸~mT#��̂��������CN��C�D��� %lǸO@� 73,��6��y���Z�jzx*��9��ʀJ�����2�0�|"AE�˸�+5^��-����r'�ۗG��o������ z�n�cc+	|cR$	�ap�LU����˥8�C��V?��>��e�@4�Ƃԁ��x�S�e�	VC�(�<X4����|/�ID����8h��AN0���4�8h,YH��1�kJ���'�;�{�J��c{)&��|��7�^�e��3+�NA��xw(:�_�л�ˡY�<���**�q��`1/��~��LUY�]����&�ϒԤ���ܮ�1�a;�AƦ0!3����JP�㛙�6�2с�lL��'CC�b�o+��q��3gNW��������[��Eco3M�^6ѥ*���K�D�X�s^���=ҷ��p�	B9��Փy��ԏ���x7jq�r�>�B��߬��!#�}��g�]���������%�}�#�wԺ2SG?��/�:#�D7��D���ػ�1���Ȱ?(��t\>����a�w�T/Q|L��"}w-��t� �?��114�ƫݚ��,�യF�gm�M���V�� #-K1�,Mejw鋨��eǕ{ݣu�c77n��.f���`'�#�ϐ=##�Z�/������D�7qq��E��W����+Աb���q&�:�kI8�f}�*r��l�p}Չ�8���/>�w�w� עV~���і��/�qz�V�����
ea^�V<�S'9&�vB�tTd��A-"�^���hS�t�t>�YY���MBC�[2{�i�a���BѮ��V@�r�PN���#�ʎ�p�,ݿ+Ϊ�*v;8Cp*�k��Һ��AWF���h�0��+�'m� Ze+I^�E��[Έ�jߦ�(p�C��~n��eĶ���%3��;��F�xM>;Ώ#�S8I_B��R���m3�������|z?��OA�>I.*,|���?��n��0-3, �,�����`��g���Ն���5+��C]�צ{�6C�&DU�J1ͼ��^�)g�����Xy�������/>0�Y�Q�ִdi��8�H�2�hd�&�d݉�:�wPY���k$R��\&Z�Ϝ7͉F�2��Q1�pӲ/�!|1���Y�*R��/{M�H۴�� !���4c�"��D�/ZF-�5�C�+G���c� ������R�.ť�Q�zQ�)���41l�<�$Qm�k�ݧ��8��p���.i?]�+�cձ�s�Wd\p.Y� �"�2����\tw�5#Ƽ��Å�z���l�W.�l*e�����8cD4�<�~���>��k8bV^m.7~8b(�������i�!�7�*y�O���2�7 �.��vl�k�t�:�j��Μb� ��eas�l�<�@x�|�&��o+o��� ���Չ��5��|�)g��8�&��� EC>5�᱌�j�֍^���|��k E�Y�o�� l�L����ĺ<�0� �WOc0	ߵl"jgK������>"K��Ly��y&�B��
m6��݂b���2Ø�}r�h=Tt���C�,��!�g8�he���ow!��BY�D
��y\����淁ڐ��$_���c=�aE�X?�}���-�ȴUK�0#�����E�lvP�ߍ�̰	����VECLh��?߃~�Z	\�A[��R�x1F���ӄ-�êC����K^$�
���I7�m�"2��kx�!�����Lt�u�T�$���63�f�7�flv�X�t��r�}vk�K�rZ���J���)�Stt9�e#(GdQo3��Y̴q[TX�)�]���=����(A�	�a$5b��z�<'��祴CI���5D��f4x��'O+�:%�t�FS<L��cŔE����s� 6�v�����Q�Y�w\m��)�
i�I�p�Mzh\�!�1�����=c��B�{3�����d�D�ԁ�U�q���&d&=�^����#��o�\���Rm����pN�c��&��ct�h��9� �U���]�7&����$���×�~nؙQ�|I�����6`Kг��W� n��6pl�!�1)أ�up"��{�7Ea��T�Q6xd�=��e����ۀ����ḋ�\����T�K+�e����v��f��D|9�:Q�	�j���Ǭ"���Ptvb1�W��gp��Ԓ�M`}#�{�g~:Sٙ����������|ұ�$�zQ3;��ݦ�<u_`�V���%��d���UA�D�p�=�筟���gȢ2 �N���5���Ҷ�ڮ��`&�$z�)�*���)�!�Lu3�G�i�=n��}�E�C�A	gtc�T����p�P��ã�)&> ��Â����ҵ�?etR*�4m��#�{9��9n������J7�� �\J��R�;����U
@~�b^0�bB����͢V��k�����7�r0X �ߔ���|G��H�8�����e2i��-�OZ������ތ6)��A!F�,;�[Ӳlp��F�u;��\<E�jXV�=�t�`�n2I9%�S�\��� ���W@aD�=��\�����+��	�zH�K��Lf�Eɓn�M����1�\��X��V���	�>WX�kg�!.�I-r��9�%�f͇�[:jak��i��[�+���4�؉Ȑ���[k6*�8�ɶ�"�����q.p�O;����!}si"/M��pW`���j�R�r�}}�U��O D.}aV�����1\���{d�ϗ�.�YZ��j��u�F�~�h���#�l$�����~X�U��V�5��w潽�#�,K���b_\���t���H��\��Ry�����E��P�_�<�9��@e�j�7���+T��>���X[��`�T���V8h>4�
�$9vE?��#�����4 ��9O4'�:Ƹ~:f�ȓi�r��6GG�!�d�v�8�X~�Q���Ը��eG2��_�,���4�~KU�d�e�s�2�X��8�)7WY����KmbPX���ps;
 K+���a�n�����e�|8i<�1���$�D-�����}�:�J ���J�
c��\���q�vEG	�E��	+1�1�|7/��T	y=.e-ܸ`W	���dP��1��s��� wL�_7�~�f�~YO�遧��c<c��NX���s��x� %��`�m4Cs[zbTS���A�Q{����Pp "J�~ښ5:�sq�}	*����h�R�����@y�2�,1yM�5���}{�i�ʴ�a)
=c�e�%�u�	`�|'P���u���e
�����Ş��^�̆�Q��x�;7�Ϛ�4�JFӟ��\���ՍY�Y[�Er���^��?��5au�'�5X�Y��i�G��כ�ڣ���{^��(;��R j;1�nz."�툏bf0�;�1�����XJ0�u�+�ҳF��]4�_���c�x@��7���d㡆�BN��T+������N�U��6�s��_Z,�Hg�T�hUw:;X�4�Ga,��܍=$N��oߥ7~
��Z7�}�Kh(a�I�����V?�M"_��T��?�R��v<����>�B=(�M�8߆!l�x�Ϻ�P�������Hւ?���Gz�aC�<�KR�m�� �yM~l��9h������!c@��67�IRh���>�n��y���V���UB��x_��V��s�Nk��]���� �!�_FT9��L��`h���B@2�9�U+?���a<��.#	!���U�ѓ���՘����:�[$)>~$�<Ɋ�8 �S�cr���z�$�L&���2���y�zזb8D�0F��f13ؘ�e��q��𥵾���\�!��%�=�6�#A�������4D�<o9�x<#���V��d�N$]v��T��R5�薯)z�}�9)/��Ќ+��*��ˆ�S����&�j���鞽���Q��ƋQ��KJp2�^�!�-��Eߢ��꥓}Z��6V�'z�PAE~��į�ʟm�t|V3Π�)�޶XQ^���M��!�}x�`�`���|��y	B��d�~9��F3r� ���.�r3Ty3K57��g����_�z�fV_`��!Z�����w�k����u�@��Iƭi�l{�8���G*��\��&�1��Ȁ�P�V��}*��,�/�`bn�ZW��~t�o�~1gg{�R_���G3\���c��C�����B�#�'�ˬ��%��Ó�fϩ�j�̶�`�,i�TQ}1Nh��+��:+>fk��v�C uY�?a^Ԧ���]o|�\׬��ZI$�
��<�a_n�� }^q��Z�?z��ʢr�BGH_�y��l����ڵQh�iZ%��r��n�gh�<Q�����s����I�0��Y��;n�U���"�V��J�c��;}�E�(~0>�r\BL���.}|í���dD�2M�WmXD���8q��D�8Ĳ��e�#�h^��]	���(?���i��9���:�b]�b��F%�C�e�����oR���!�!�K��(Bۻ{"��_;nKyli܆py�������Ȉ�}�ex�#�-��W�٫N�	d�ss�bf�QFQ�E���\Y�ڐȀ�Q��JZ��c�V�
+(���q�Y�/UF{��K,t�b�N���4``�}�*o-��_c�0a��,n��>?�O��F�EH���������g��b_�OHGڻ�so�6�7B�/�J\�Y?*��]Zh��^�a���Z���<^H��ŭL��e���롞��¬KAL��V�mM%x����݌���� r|���C&�����(���M; {I����E��#q�n5įD�I*z�O��~�?�7,��OɅ�dDǝK����	Kh��ZG��w�1���X)p��?a֦�����%P$��D�_� .>�n�en$G	�w��cB�G��3Pr8���g4:Tk�65�Za���Zm�x�#�����d��6�ۋҕ�deO�͆/�����Ě�b����/C�eq��kA4�bd"߶����S�^z��>f�Y���+�AV�h��n����Q��*�
ˋ?m�<�1�@��s���q��:��dP�(���gB��.����U��a�6}�r����v�X����>��
&���|���@|jq�q�R��OKǅ�W�-���1�"bC\�R��sQ���%&��B~�Q������w����A�ʲg��T(oS�8:&�N��p���:\U����cŭ��q�	���>��X�޹��y~�0O�5�����Fk��ρ���T@7R�<jd���KJ�w��%&sOwe%�g� ���^X��=tiK��Ͽ	#X�ʞO��*547򺅘��~��?�#��H�?3�n����[�]�w3�^l;�%��#isE�c{��v�t[x.�'���0X�t�H"A�D�5u<��G�) _���S���}��n���l���; �;�*����_�bd$�U������L|��t���*K��%�Bbt�����S�i�F��Kn��51�	P�W���C�<�X�'4�2��e�H��%7`g N/�t@lF�X%��ŵ���B�:Ȫ>z�|�m��͢}},�~	��].�YWl�+�n�.�v�36��)���B���ƫ[5ȵ�M�~b�}���խ��|�X�� w>����*�4�d�Pt�,q|܃��؝>�Zr��	���?`����p �:=�.��D�7�\����.h^���dW�dX|����jM?A�:��>K�m�g'�,�IzV-El[ef�j�*���JJv����[���[:��%��|���*,�p<�+�?5���EVt-�Ѩo@2F8!��e`�ׂ��&���l�P�#$a|Q����=��ޡZ�Q��Ly��ˎ�+p��pJb�p�T��ϯ�(c[����pE[��qV���7��Q���x9���@I��|�l-}�+�b¹�2��ރ��J��w����d[��d�4�b� �H;:���9�,4L�Ed���t���������2�?�'h#+Ou�a���1`~��r-��cF�gƍ�WO�f�%��\��eK�Z�(
�v�'�G��}U	��q��2���uM���v�a$��`Lm׏���l���4Q�W�9!$��S7�@�Y���|5�=�DX�]mI=��J�C+є*`���	�a���`BWO&5����ւ9q���Oj�s�\T��C��3^�d�����_��xJ���3Z B,#x���酩K�g��m��=��j��w�z�y`��Ln�,l��f?N6+�c�%E��F�s��� >�Q�σ�L��_I��(�������	`e ~���t{ic��ʸ��⫎/No^n�^�L~4�F@��5{�m"q���._cX���,*�t���&�{�+��V�ܕ��>�|�R�l��Y�_{n&K�h�W�]0��V%~=�z�K�t |�*Դ#�h�ᴌ�Kf��T�Hw��Fdg�Ԯ��Y-�_|�$������1����쥌X��:w������\�0?����r`:�wl93x�.v�ml�N�F���b�i�E�R��z�ML?��ĉ�fâ��"�'��Yt��{	��h�X�1�o�cUđ�x3��#���GA�7R�B�=њ1�7���ԁ@���	����vo-��
7��O��N����1r���IG�Z]g߆r�aq��.5�jw�
+�՚>Җ�Q��j��*F�Y'0Fo.ҕ���R��!�)��B @�N��H�'>����.XH�4G���	�^��P[���W ��N�?�@���z�{�Q����Mk2��]�ߚ+��x��N��$�&��C�mj`br7��E��`�E[kDT�����%�XϩY�m ��-�;pe1y"�p�e��^zi6c����D��,kr����t8@��9�C��ϨLI��LCH��~�`zTƨ.F��}���ч�X���6�[g�A���V�����mJؓ75�Z�ƺ�0_[�.������iq,\y�W��u_��Ĳ�lOz��xjO�����k|�8>!�5�����r.
�����{c�ȪO�9'I��p�����p�Hx���@��Q�f���]��������Al��
4�Ca�^�.)k�y�!��}(ޮOJ���̱�+rd���-q�_�j���ҪI�q�O2Y��ƉB��H�`z��0:���a�W�Ɔ�\�J6&!=m���IE{��!���ߙ�ڠ�H̙�����G+c0���l��^�~�Н����s>CT��p�J]��ҵV��A�*x�����;�������]y}�M$�q^�UU��:و�ҏ�
�t;�'�t�@�����I�7��iP>�L��+;�7p�>��4�F�0<��ls@(L�j��ߴ��i�Ak|��q/J�W�CǾ��!擄�����b�vV��<�xA�B>k�q�M9,�M=��ZφTSB��.}3o��$�2)#bJ�$��k��4b���?[���^E���I�7��-ۓ�0Z%�[)V�S
'v��Y��?�B�;��u,^v�ᕴ�����y&������Ej����Wh ij3�B�a��#�LY��A1?�UN�{���z���R���8yG�uR�����7�@ʭ���j��I����Z��ݖ�u��n,��*��,n%�|�ɿ%���V���S2�����^-鴣�;dr�-�;A�S/;�x��\�Lf �$�|�բ1>� ��>W��Vx֬ޥ�I�;a���6^���rq�I�B�-c1�Z0HJ M"�2�P�힖���G�����C cCm�%{L�ӻ�m�n�gY.@ݳo�pV�����0�;����V��9�T"���KUJ��i�@�*����l�����`h��Ē���S���n�]�����M��E	"[�;����΋���~�̘H�B,��I0�v?����7bN��e���)|I�ʤ�����2�23s�й����I���Ս�GI�g�N�f��'QBf���������p�>C��=�{�Wi<���*�kT�:�z�?���^��D���sdo����*x	�E,7���"�\[TL�_.�([�SK���j��9���Ȓ��A�8�+[��.�$�W�d���V��"C)���5ESN�>�PN<�#?�|]y"�ן���=��LNC�������hM뮺��ĝ9��1L

���81М��b�d��W���og�p(�A4�2�"歇�Lf��}�*J矎;�����2����G\k/���y�-b�60{I����VL[V�y)���_�x[�
��ՇIbI�V�l��w�K��^t����fX�k�Sv���y�����ᓵ1]s��!9����uEI�V�W�� ���&`�{�w0�"8�`�'LW)�?���J�`�lƦ᭤���0x �kz��-+�����+�]%d��&�!�3���O��Ǯ�����>;�N�@��Ծ�ЗA�_u���A9t*���%a��0h�M�e-����+�]I�V����Q�1���۸�|�
S���7h�S%�0B��;��z��b��5,�;���A�+H�?3�n-K܏'�9�,�k�0���v�$W�M
x&�ԟY�L�T��>*d���l/�����%1��hFv�=M�=��T�<��3�|�ia�U�������j�O�y'���dWpcGl2Z��oк|ɢ���7�v۬(©��Ɩ �A]�a�	�-$
�Y����L��h"N��XZ�q�-tj�,D�mf6{VQ�cr�.H�zZ�A��<A��z	�F���oH��̩��c~h��,�>5P�%�P���=�XX~�?�1[�߮�T�O�ޡKw!��c1#6�a�@A|��6ܧ�<�c4�zU��@U�N�@�'T���osn�%�wE�\��}�vf�Ӌј����� �A?d`Q�����l�8qcҗ���_::! W�66���8���#*ǫ�WS��Yj��i��j��pṘ#�t�S@���$l,,�b�g�-q��3)dk�A4�gA�fw���f!A��Pʐk�}j>�'�E��<���
+ox������{�vF.l�c	�E�pvq��3}P`]Y����{���r�7��b�3�ɠ|Gs�}&d���Za�	HzOf�P$}^s�-Z4A��n�t��U �|�
�yT�i��"d�0
��uE�]�
�m�D����D\a��`O�ʝ�V�B��Q��"�����ڷ~�V��ϣz��a�;q^� ��Zn�r7�����0���l6��a��p�e�Ʋ�C�����X��o{z����ܤ�0���dI�v�Ո������INO���3j���=S�=�h,r��6p��-��*�d��m�r�(�ͳ�	$�˳�=��xV8��h����-��+ǫhi�f��H_�5|���������&��v�\jo��Z�0=#73�
��$���k ��G�޲K�p�6?-O�ׇ$n��1���e��Ww�9)�׬
-SCѓ=��JװCn�~��h��}��dw
���8GGbd��d�������pC�t,�!7I��+
�������0��`�IV(� �Pǎ�:��h����'�~M���R�D��ls��@����u�ON����v!����s�/x<��������	8�}pf�l_�ؘ.u��lHXx#f~�)ydef�:���d������̐`�pnA�DI�/~s:���R��m�cc����#Vce�D,BC������y9�Id�� ��� �Hs����In��luS��&+����@�p��KC^W�O�Xtlݰ���D��-9	h2��(�v[�d �(Qjn_b��>X����H�
��.o6(h�0���$s��o��#��e��p$�ΐ��wHʯ���6S�P�,d��T(m>���-1���`�~�
P߇���I�<[�<�4%�J��t#�,�� y���m����G:�@c���uK���H*f��w���V���t�?J���<�,N�9��j��V�ӄ���F�j��tM7/�XbYҊXX�jh��B۳Pcq֞���������V�abLnM7!�k�t�����G@�Ruo*��T��ww�:V�1�,{� ��� *C�Vce�5ʟ��c�
eU�¥����4%�G��n��=NP��^� ��� 	� $l)�:De)���	�Y�<������'���g��]���ÿ�06n�>�l�Ȥ;�<��8���]�Jt#\Ȍ�9\�?LH �+��jl++�V�l�52&+������?�/s��F,1�J������Կ����2aC���O�ɻ�T%�����in�_]B�a���b�3 6OHw>b
Է����CO�˾+�����,P).38���y6<�T�[D΍���)�I�ت�P����:'ƨS�)��?�p/�e���L����������]z��w�ְMVM��~;��p�� $a�%��|�3�L�d�ʼ�~�e�'1)ī�n�K��g�قX[t����¹�cfǣe�MѪ�e�J�`���c7�ݢ��,ԗ�q�����QI��uǵ�؈h�sF�U�XT�ȕ�Δ�k�}�z�v�T-�hGP�gq8� �r���Wu��C�*�)���=��[��tݶ�PS@�A�U����!Y��6qec��^K[�ß�xhFդUV9�7���ڐx�F��]�:�: n��8��Z���:t�ؑk�.?ӅP����W/>$ٗ������uh��������T�c'`�G������.?��|0?�@5?<��G�޳�1��|}����p�c���|�QBڧ=	�����k~|촅T��B�[��6g+��ːC��jlKXRwک�{�?��e�_���U� 0]�݊���4S:r�_��e�74*��@��,m�/�,E�|����
��
�m�|9�aY>D��"�]�b"�hx�P�R�_jN����a~<��xK���v��^e�u*V���@R���9�b3���:�j��Ѡ�5j�&�Q������dL��t&ٺ��:�����Y�F�Y����?�&�s0j��Ȋ��G�L�7>�������	������f"��ĕbZ�Q֨�6k^�����$��=�V�<Rt�&-�wg�2?���Q����j�q���uPEP�P�	�Y�E����d���:_M�����<bD���T�{�ì|`/d�pj�pS�n�8�%\c`��܃�DK�S�8{�h�6��;CR�������+��l��ELbf(�0���M1�>�l�N��Ȋ�V���@u�y�U��i�G�J��m.!��s��@�V���I,�s����w�R1&��wf��O���"���H(�������_�i�˼7l����E9�-@�7���jv�#���m �K9ݞpkVv �K(J���%�$�$�������|f��Uy�a��F�5+�L�?�aKh�*>���v��DO��쬱������8a�뛙9Y4�~��m,|^�#���u�*l\����udN.�vl:�}h����?s�9������<���#����^MG�L�9�l�V�4/3���6�� �ϙXx���z�ȕ�Mk3/�	KcJ�Чs�B,��;�)�s�"Z�	���v�m)�B�D �Ǟ�,^�����2�&^>z�H�2Y?؛RJs�1����5�%�D�!F�$�"����<���Ռ<��=�� ��9���.�JOG�H�F�(�,��k��q�TF�dz�Ԍ���w����F�g��x_1+,\����!��0nv&�i�%�� ��-n�o.�h�H*׮6��g�~�7פ���[Q����`�7K�E��/�ȑ��=�n0��T��5 êtL�#���:|~��GPz��s��܈���)6���)o8֢U���P<�i���v^�r�?��'�@�/Vk�,�q�	*1��oX�z))'����ZTf	�S���C����6��1X�\�;&Al^�-g�#>'�XO�>���P��n>����O�:Ӄ���?/*q��ِ�� N��� �H��jR@B/�^R��;'P�^a?�/��3ac�1�������dǎU�?���[�}�
G�o�c��v����Nj��Xl�_a���W�-޹������1�����g�//#���D�>����oqBޯa��LE����8���=c�����zҘk�kaV�9��G��QC'����_ sTL����O�(�<��:j�K�:Cɐ� ���@�1NV�u᫁� t<���YiF�QM��ҹn*w�9T��M�o�hq��t���S��_oOD���B
ݰuc.}��JT,�<yd�d�YJ�4���l���y��)%u.��"|�
�����7���{E���g?z��X`K��q]�����$om�UE��0)��R~�X<3:�
19y��A�9?^�lG�M>3�J�ʠ�_���j2�U
�/h�� �K[�ƿ�C?��\�T1���(��i{
?o٣/~ �	*��+W��z��vYg,O(�i�� �:�bu|)\�E5��S���������Dh� �F-YxRX��_DW�s���׶�`p4{r��ިb���
<v�<c|� {ĪL��i��
�Bլ2���w��!�X%�Կ�V�Q��~�>�+SKH�0�'�s`{Hד� Z�<x����F�Ｍ�d6��*��<}V��i�M�H=���j=w����@�o�T�셛>������+��ƽ�9���&AS�a����7Дu���v-�����n���]��ocBЛm�ºPv�E�6)=�z����L����S̂��KE���.�"x�y�Y�_�=c��jk�B��7�@�
��5q�ehOy���@���ܼA�z��AȜbQ�*A��g��&/�a�����em�V/�����AT;e-�h��,g%d����D�h�z.ޛ����l�D�����a�LI�V�ѴE��l��`�ꁤQ�/$���վ3�Lv��>�J��6}jʃkU�֏y�~�|=c���I���\�f^mbM&���m`�cXG3���p I���x>Ubϱ>	���<��S���"�ٹ����F�yR*�����F�K3b�@B�t{��ʀ\���͐�N�lt$[�H����2	��t1����e~x��[�b'���n/�ſ���͘I�&PS�N���q�o��PĆ��>s/���f�'���I��' =��`�E�S�#Ͷ,k8H��X�S�V���P�@-�;�i��]><#]PaP�o�J���^9�~9x�ݽgq3D2���Cˆ��ް��H���9ķ.b� .�01h��@� ��&�$tÝ&��;�h:�l�����/�!%�K
07���-��qA�+ҥ$_x��潾�@�J������
t;�0~��0,�Ñ�֌D��)V����x|��:|�wz��￰1��5�����FmENl�������ml��:
����ЯM]�r���գn����X��7�nj]?�k�| 
\��vl~���e��Jsb��7C�a4��O
�Q�~4�Yh>��)��R;�*���,�1������B�=YЙ��K(
2�<[,�ll-���FF�h8��&rl�搨���CY ����GY���M�63Sڽ�I�ةX5�W�F ��&A�v�>�9䋓
��Ǭ?���?����	ʉ#�Gk��(K'�Y�?�IǓ��!&�5u�.y7>OG�]'~'��+�Ձܛ�{�Hq����z������W���g�u%��je\��U��kh �_��$�f��I��Y(�'��i���uE��#��oa'��S9�~(��E��c������fO��������E�V�+�Fj������A6l���Q�������� �K��#�Z��"��ح+/lL�X��4tʴ�*�� *b3� 7\�I�2���J/��_-g��7^N�r�֠�2��f4 Ib���`�ѕca�o��5cԣ������һ��nJyኜ|Ш���~��ГQ{l��N&(/���(�pMB��㜯��6��@=���5�a���{���l|pƑGO��J��C����n-
�!��ѭ��BrH͖-`�{Y�����J̹��e��vy�!����o�ߒv[�̇B�X=���Z'L)�����Y�v�sY]*�q)-�o��������� ��a�v���<.<H��o@�x�5|+Aqj��e5U��-�K#),mU8�K``Q�{C�-_�x�W}��_��=���9ϧ���q=��'��ц����ft�D�k��B�Z��6���ș�發!�O�/e��[��4�������-�x�gz6�y��uJ0Ѧ1����?��Z��k�g~m�c%e��� �b��%���"�o������l㥌Q�I%���8%	�͐DG(���Z�G��7ң3F�0��y��}��i�Ji�_�db��^o�]|m����ƺ��Ҍ#��Y�	�����E�|}m�ND�!U���o[Dҧu_��Wgpʾ��K�1$��v�R�$֘:d!s����b|�NǦ,V*նl���V�A�W.���S�� �%�K�x�p��lD�c�(�O��B���Me))�"cO�J(�'�.�@y����U��v^�}���:S)���u����f��(#����8�ɇC�s=�fr�?N5M����Ia�(#*U%P]h��ُ52�DAH�c�IUr�'X�2��Qܧ�z��ب"l~�i[t��Vrc� �ba��*%�U�$�J&w��0�1=)o�_�ˆ�ֽ�߁��s���u����&f���CI���'PμvƊ/o�r�'��`nb�lE�ʹ�_{-ƍ5�Ӆ|F�EZ���m���T��� ����"��O��V��LnIw�{Ѩ��X����W7�|X`a���Uņ��u�9Ι��¾-�_3LM�	����(��֒x����^=�i$^�j�bP���⟂6��MK�����t�)��M>W�XED�|�ݠ/�Q����͑,x:L���,�^r�=N�q�M/=J�p�D�
�UB�
E��[bS�Bj�	�Y�~�	5hM
AR��lRn�$�q��RD6<�D�~����r��Ax��lmc3t ��OWf�^`��u��~$��Ȍ�g&�{���R4����	U�[#��u�2i3%W�09�E��w�h�xg��^�џ�<xw��m���K*�0��74k@Z��if�`�n�9?TMK��9I������4�H�� �`�����U^ʙ�S���ĄJ��~�=n��	g�jnk�;_��J4it;F/���'��h�ԧڞ���4ߠ~'�4��H@�0���|� � :��/Ӝ�&\z#���Lr�;]�Zq��-�!L�UN4ba�D���jr�LB�}���
�q+�߮�?L�t�Q_[�A���K�U��U;@C��>�L|	�?g�*��d�)���d�%���Ʈ&��&"�z���ۦW��Y����[�шI�x��$��0
Cz��������MԪ�����)7%R%܋��X_\kX�f�]D��N��W#�(E�H��ٯ���ygT�$u�w�|��؃�D[��?�)�ײ{���e�Z&Om9;ٴ'����"9���̖s�~����7�?����)M���'���bCbL}g���'�`��̧N�U�B�&�b���>XWu<��MQ��rIw8;�JI,R�Z�Q��ڱw��O[�g� ��b��*ƭ�%D+���]}fp�&\?Vf��1W��l$���]�%��'2Z�Z�[D�x��(2��x��5�j�K�R rm��5���Ə/|���@r�w�;�(#q��z7�ZrL�	�Ɗ/W|Sd��C/�Nuɝ�	ʪA&+�4x��<	sv�~9~��Ӽ�+g�1��5��i|�Yۅ�c�y�H^�4&}�R��1~ �ެ"F~:y/��̲���6;ud�aIt�Ӳs3�j �`����G��8T6�e�Xnk��g�cc�ȥeS#��M����K^��;+ۨ5
�z��XC�j��O[x���]��ս��껕<�'H\�ܤ�@}-]-}�����'��f�;`)
}����$W����-��F�hN��7>Z��-嘲�㡑I�r��V�;�F�ř&���
W�<dL�Ka/�Pv"�u���IW�O{���+����i|�ӓ�ѩ�"��u���0Lmwl���c�'����3>F�x����?��t���J��áT��e���|��n>�_�U�@_����#8e�
У�WQ���,���bn3G\}p��\��{��a�D�$�H�CV�xּin]�H`P���348�
��3.�!�ۍ���z�`��`a+s����aF�G��O����u�$��l�`S���:+F�r@�?�����ْheC��
X{����k�ޗ4<�Y���u��ׇ��A���D\L�� �X���n�?�-g�j�z�}���In�#�Wp]"����f�J{P�^Du'��^&���g]�B��G�v�ɅA P	K��R�w�%���?��b�j3K��5�D
R�@�F�1�b��'Rxg��g	����I����*�

`%�(��r
p���(�*Z%.�`�����{�CPH�](�����T�-Y\�Y����2�,��)�?�H�@������)�"�D�æW��ܕ�D,ji��Д�G���{��P�'�Vt߭Y	Yts)��!Iet���K�a�=aK�H�Q���Uv�]��o _�L�+E���a?��ڇ�`���4-fX�?8�~�<
AHO���c�_=�A�B�З�l�''���-�RE[?�2o���!a��##�l��\��Gm6���y\A�V��ި
+����+!�v�Gu�������ο�s��yoB,WO��KN����{�X�ΐ(C��}��y�cq���<�ͭ<�
6�z�(y��m���]%�:*oW��1��M*��MWY����H�l<�ˌ%-׮�4\[�tɯ�G�=�Q��[��R����@0���W��<x�E�N�\T�������1�α��"
�?id+����ˢ	�{q��/�V �-�E��LC�R�.�q8����8�/�Vn�?�9XCh���;ץ��d^�J(ޱ�M0Vbe8��5U����%���/���n?��Ϡ�
:T�4ջ�@N����F�f2� Sq��O��B4�_��{��#��e�|�K��3 �Rc��U4z��pdQ�NNإG��:��DT��ݶ��g縳ɞ`v�.{@El�U��)��]ۣ�1�_��})��g��V�:��E��%���h\H�ɢ��~��H�)���w�H���dh�Jo��Y���9<�fS�N̋D�/c�k6M~ê�^9ە�8��9SU7q0�w�2~ "��t��c���(&$�&�ѪG	��8�j�7H�_(��v\tc�4���������h��1��A`�X�C��ѷ5O���w �-Ų骪�^hrn��ˡ�x��%Ϟ������=%г���S���aN)g#�|0�
�x\��3]�f��3ن�\E[�Eg��egM*�z��k����Ǚ��T ,gKS*��ߚ��u2ڵ�I�pL�!��?B�F�uz9�s(�]����9+�H~��m!����?�\�=����vK���|�@NH�� ��y@�*��{�����˺lQ�m�rp$��B��U��E>u��@P��N��׾;D��^$���g{��f�:�@;�,�ao2j�=�)#�Lo��tbe���}.-��0�0b�B'&�H꽰������T�'���f-����$���1�����Z䢝��Y�U�&��|˽m'?I�?�*L,h��)��|���0݌���� ��m�"#���,�?c"'fV�h�|��q>9u#�Ψ����Q���s�4�.�A�a���|lG�	�(�5Iwƭ��NnM�9~d�?��DQ%n�4*.Pz���	|���6��P�q�jx;�^�y�/{\ O|<.�K��V�}R��[�v���!�TM#�j\(GiMM7�|��}���+�5KWV �Q&�{!�/�ͨ���E���	$c<��A�������ȵ&�M{⻰��g�Dn'�u��$�jK��̗Ε�7Я��U��4čkmvP��ã��A�[9꺃��6���19��������x�M�0�#�� �DȘ˛���9�*s�̺4��G�Wc>)n�8`����P9*�ZF*�*}B�ȯ5��>o� �� JC/豷���G�r�"lμ�w��<�"2 @�$�h����z�Ԥ�r�A�����vV�x�:"��'I�zf�m�{	<x�A=`eBh;���vGol��J';���Ͱ��z�Y�'�zJ1�/�2��+!,�g��.�@��|�P���¦I.�t�����xo�?�[������f�M��E�t�(�������=��C�Y���7L���Q0��sڗL�y04"�{��d���^���.��R�z����Ns�!�F�a��X����J���Ц��g�<>���^�V)�ҹ^�,��U���+�X�X��ߤ��e���r���ā7W�K��b|fٷ�ˮ��K��f�����9�&LzC�3�oL��ߒy��{�	�q9��%��V��^̤���Y�����t��g���183\�9BS&��M�(�_�"f�3�ي�aW���<��,��EK�����[��Yz~+	�-�R��] R{׏��)����B(eyT�˼n!����� �R�؟&[��0"�c!��)��i�+1�5���+f�f�(��~����yj��O��[���ǲ�RL�nZ�,(��uk�Z�nܔ�ĭ�0��N���4Ym�t=�C,T��~{��Cf�ۭ��K�����H��_�4L�3�=��u��
å���e�;�_�r��7-�t4h�q� �sN{ʎz�|zK�%�$����?�~�c��j�r�ڏ.2�"�sS�G�I��z0�E'�D��
֔�6j�Qy��tp��(����&�^:����?��K��@,Q�j�Yіi��a��[P���������[3���%�F�� ���eR�3�˩2�)N��]�O^�b�r��s��k	ŁH;�]�!���7I��]c�����s:�u��Y��B{.�Z濉\��P��bz�iP���I����,ltP����ЁGE�(�v]j�Ƞ��r��'/YU�XO������ �(,���B�6zK�l&m�$������M�e�,�,W		���E/QOJ"b6�Ҳ��[�ap�ѭ�D�:�7ݕ�Kb%�������������y���.��cu���j��"��Q�Nq�=�`�A&���CI* ���� ��8|���W�]5����w �����x`'w�@�����KH
�cb���s�ȫSɿ�4�5�s���")������pU�lf�7Ȥ�N���`Z�p��GA���U�ׂ���"t�B��,�
�-���u��ٴ�>�2#�n`��.�����&S�T5����(�,��.WTO�m�\Q��F�i���..���vw�v!�QVoA��FTM�e��ǽD2a�"ꀁ&��2#�Q��
:p�qA���&<�6��������^_�Y1���h�!#}]��˝��_�e�>n��o4V���2��,�}9�ni\�d��/39�i���Z�e�q,��͐�|P��� �������%��3*�W�5�?�C�O�B��m�Ul��[�!�������\m�V���(�
����i6�N��K2Wп �$�����'��IP�q�\�?�Jx&���d�o�EW�[�~� R�-U�� ��68�a�����Eޭ���UkN�ud�{�hetp��!�e�-
;l7+՚�Ϩ ����6��04ɍ��֓_��Ҟ=�U�L*�D/U�֑5g����W�m�wut�֮�7/(��7�9�G7�SZ2�2.������=a|���"��\�7�~��%��V�����G�_"�{�A�K��V@�)r�}�o�>�h�P&Dv�s.�4�%1��ޘ\'u�xi*ίN��6���2��o�9�瑝g�vȬ k�Gp�����Q��s�O���%&�(�P��7?JdF��1��΃+"!&䪂y��<~�Љ[�c�,Yh�h;Ѣ��0������U�`ؐ�bφ��1�|���SyI� �z���U�܉.j��V���)R��7x���lر}��������~���ݞ3]@�tH�+$U�
-"=�-(�(������<�Я\E>=fF<x�W�����ӷ�:���
S�&��.��_fg��q /���ЁVl!�,lxL_��fi��n�ǘ����'8렻����mr�EI��b�\����	��c�ͺ�k<g+{f�`�eo��J?� >�kƁ4!i_�ƭ��vG�j�:$z��+<�Z�ȅO_3��'s���3xD�ڲx���~���"d���F�=�>g���R�3��b �G�)����]�0u�'~����B祮q��3����WUQ{����@�q M7v:�kY������ws�
�sz��Mt$�Xi�s���C�&�}��K�e��c�/�ĵ��=MK������#��ņ�0�%�É��`�R�1A8��f�HQni`��P-�j�<���g�63��6���s0G$�UM@Kl|y_�`iT�Y�়�4�ύT�@��0�����%���ER?p\&(�� y+|����]㇀Dz�\�ܦz��=М
���zEư�Y���>y��-4�ě�sՉ�rA��+��2�ħ���x���� /�
L��̓��"I���㒦��3>���Q���4n�E��S~�w�t�����N���u��e�0~��D
ɹeæ��4OǇ�q@OVmr`���"��ߩ��t+񰹝�s�� �n�Y� �L�@t�\�T�1,}�z;�9�(��3 �B��Ѽ���|��T%T�*0.r"9'U�#ˊW]MK���n���n�ܠ�]��1Ѩ�m:S�����8���5Qg�}!^�EUи'L@�x$��g/�`���=����EA�	gG�:#������|?��_]���aT@��Ic6"L\��]��s,� h'�պ�g�G��r�����MWIF�����9�6����\W0*Y\�ݶ��3�!*!�:�E�R<+�%:����a�Z3��#��-���%} ���v
P�J�.2��t�ϛ�H�v�~��qM$� ��`�*���)�^M1}��6�{ �[�3�f7��� W�'O�q�j��,鬫\1n}�z�@~����z��������	�[X��^c�vx5(�uP�n�<zK���!�<>��)d[:���`�
�<�2�2�9����c�H�\��I����jS+�q�8�w�I!���D8��5�7���h���G���,oc̬)��@�����x���#���ȬtD�Ex������[v�RV��aB�$>"gQi��\{,#�H�Պ�Ų��ˍ�
F�K҉W�F�m0|��ߵc�:rK]_nY�Q�93`�It&�ר���L���I��%�LU
�8SM�⭮�8�؋�hT]����8�'C�#�QX�<'mT�Kq5�L���М��������������R/ezOX�T׎m�[�2ܫ�X�T� έ��ҸB�R���&u?T�"I�6|;�?�ƅ�N_��o��؎q&\S�e����W�w���cQyL��$Zn�`K��5�6/�
s��M����TJ(���8' tՄ���/�����n'�X��e$ۉ�<{*WZ\�~�F��<���}�ow
V~�9㫧4��d��{ U�q��Sj��d-eʄ.�0U?m��1��$Iu,�v��er���7�i����D�:��t���N��v*Y��-��8�IM�����d�$Ы��?rh�Z��x�s��鞨ǆ$�<$}y�ZE�*b�O��c����F���ɂPtu#�%�ڽ�ȣ-�>ʗ��C�K���[���{tݱ&��9".w8�ƙ��&ko��a�Mz~��ȭ���㞘CY�"Ӫ�HL!}�|*��H#��S��'Y_2��%�V!�����@�	<c|�/�9�U����ޱ`�s˃gg�\r>`o^�;H��a�c��sn��-:K��X^M��C#h��������$#k���EhfF���y�E�t'��"}���/��q�<��L����\�t|9�X3Xۏ�7����Y�]�;^�JS��9�\;��ʥ#wi�sa�
����X;�^�'bz>T�G��d �R�_̋n? ��M��K��ay,�E��>�n/�{�Ғ#����N`P�KV:��Έ��u��f�k��ǽU"�*�Q5��|�f�nK��X�@��;;�s���IίC�[B�Ǝ��Y�� �ߔlT��r��U^���U�Ak?*�t�%��]ŭxRH�V��4E���)?�i�𩟊2����sT:#Rr{N8-��r�UM*��wc�I�s�z�j5B�&S|��Df���^�J���HQ+U܍�G�߬�өl���Q�*q�J���s�������TY��]R{���Af���T|L�h��E���cx�0G��h.��MP^X�Wo��W@�gp����l��M~�'7�=n��e1	Ԝ��x�n+�@9��F�m{V8A��\��8C�i���-C�F���/���FBt��B�m��EY1����1�O��Kt��	��{ۻX`�W�r��Z��w�;��1�P#�b)\&���W�����{�'�'�0�ʭ�Fu�mG�X���BO�a���ȡŧ;���h�G��OM��.S�k��l���N` 娏�0�!^��p�A!c�N d��g*Z\☱U���@�o�4���;~\��-ee�e;�{�OJe�C�g�R�(O�����{��X��u
5���epj7���nZy�*¿ʜ���~�sIuM�2cұc�0�0`�b�N��'��K��g�|�Xy��i���|=��u��k�-�i�~jM��j܀�
�\	�p?���W����M����4��Bg�BA��p��۠��\i�}}���0�@������UD�}��(���:��@U����
	�� q�>�3��5I!�"�ע��v���F�<�L6@D�]�����n���)�������&��!#G�駀��ò;GzJ����Z�9�;�ݴ:�8s�+��q�y���W;�����f��f��F��/�c�r���y���5��H�xb�rZu�	��5��S"�'|~�z�܆.7�Pt���,��pׄZT�(sy����Ѽ�<�kŵ���jn'
��ĮT�կ;k%���wI/ůX�{7Q��'"���o��iQ�\[����RW�-���M��p����_����G�ݮ5Ď[�q�6r�Jf/����3�Q���Y�'��%�n��<quhg���Hm���Î�p��Ȅ�T��^w�!^�;�����K���w�W�ɩ������w������i�L����S1�H.J�wВ���y�~xس�Ã�W]�Q�=}`�#.Jz{�p��8R���1�b�CP�Ma��f+"�}l��ț�)�^�؟k�܆��g,�e�Ѽ]�	֮������3�,*@���>u1��9�E�_`q���8��n�Ŝ�����>���%>й�&������YR8�F��T���[+GS�so���Wf˺�rE�xO�2ku!��@�
7��;���-���j߾��t�di���2�uN�O��t���w������
(;�Mգm��G,^'dğ�;�zM�^y�cqبzw���E�� �d����[\�&��)�&�f.�џw�[/"���!,��~3��/a��=�n���mhx�Y����g�=F�y4��*2{�xqX�ɵ(����vR�^��E�A����Q�2p����q��Nhc�Ha�`�	ڳ�ܾ15̣������D� 
��
.>՜,��@���i|��;�d}�>BMk��V*�� o,�J��F0����D �_�����xB�7�_Ţ�~c�hJ]ƭ�����]�"�T��i�"�[D^k������q��=�YbX�Ӝ��{R���Cz��Os2 ���{��M�d�z)��4H���N�^�r8ǻǂ��d�{�O�*�|�_GM�wՖG
�o=��S��OJ��˛�G���g��Y��K<}@h��jP���9�>g�J'���a�J8�������7$N��E�d�p:������_�Y�y����\MEx�Qa���yl����p�Mm�����D� ��a��(���W<ecHcv�:���`��It,h �r�bA�Մ��s1��V�Hג��V�^�ͥf���vp��a�`�#�om��8��1(k�у^1Ȗ��4i���q��'��5�a;��m[Y��Q&G����(+������u�����PD�ܭ#e�)tmD��3Lh=Q�M���b���`E�+����-���blT��J��٦�m��C.��+p����R g�y�1�aV@��%g�BA�� � �����o�(�x�u�2|\�{����
�X;��I��gv 5�u�{9O���{= r��9�N�Kb�����C+�|5�7�YH:�x��nqn��Y>�w+�ъ��0���bR������+��N�a���g�[�]P�,�a������uSP�\X��f��f��t����Z �~�72�dN��\�3b�W���eyi4�U�3���ܱ,��{Om��f��/�����i���ŧ�-�j�O�J�������,���D;�N�xa^4̥ھ����K�@���h)d�?h���+��꫟!^�׆��ٽ6g�=Y[)�c��:�(M�Ƿ�3a�B�x�|��7��[�\&j ���<�>2�B�	3&�ź�R�p� n���js�)gCu:E����&;��Pk�g�o�!՜V#��c�wt#k�t. �(�ۖI���~L���H1b| �]��"�xȃ\Yun�qW�R�0�F翁���Мt�f�uݘ{O$���Q0�?.JZM5�V��@�h��lB���r|�[�a���"�g��������C�@�Y�jcS������*�\�ɒD���GK�k'z�6��}z4H�Gq����:T�fo$�w��)	�7��hWq��e���!}��P��J�����\"3pu{y���y��>x0b�Z8��:5��EL�^ę��`��ʈv�� ��Ǚ���>���Mi�U�0N=��L�>�մL��G���������8nN�ؿj���r�c�n�+�W�OW�p��V��p�s-��DN��_<4�w,g=�*�0��4�!��=��l

n_5XS�6j��Rp�{.2è�?d����W�]��huc�J@&��8����|�:�犯�6�U��7=�N`���>%O��!МX>�? ,����L��W�+�h�t!Zvg�����;g�NA�[�VW�G��O�����ל��r��4��. �S�v�� P�s%�w��3!���Y���xju��=0 ��L�8��@ 2L��'��"B�Nz�e��%�9�Ծg	u�l�aAQ�r���)��c��}���K�Gܰ�/v�[`o7��	=EI��}�X2��s�"��6�}{R�;�]	ӧfA�,j��sa�B�3�U�+����s�.�+�~8xA ����D�Z4O�T�Z����o�L�wp}n�GA;�\IdՑ��{~q��)��� ;uNݛ��vص>L�f6�b?��6�2ݖ0���ߕ�߾�*"Ѐ����v��<������1�Շ�a��<m�
C�����UQ�I�n�{B�#<�J��뭖T&R�]�F��b1���c0(&vp��:�![qV����\�@
{�T�����|�h<3��\�I�*�43 �$M�����,����^���1fB(|�dF����~W��0��~�)�#L(W������l|���w/�����d��.i��#���c�%<y���S����.�3�\���[#��.�'S1=Ѹ5A�����ғ�U}����	�$��?��N��P�jZ�J��� ��vC^�<��{8�clxB��T}�|p��� �K|Ց?�A����HYsc���g#�����: n���������y���uX�W��M��O��EcJ3����#�o����v� 㩎� �Fv"iKh8�i��r�Qng�=��5����P_�����l�ST2�r�Y7�	#������:�g:d�m���@ێ��jT�P��/$��e�I���=����b1��ф��wC�J�f��D�h�f�,V�ls��k��Tz`���k�i8c��|"�է0Qn���������7�~ށ�g�P	ZD���6�*���5�Ǥ��Q��dh-/h Iis��L��H숭G�l S?�x���Wv�0�a�L��=�+��iQ�P	�h���?$Y��|
]�|����
іx$�o�����4���r����:�ds�O[�c|���[�Yl�����cXN͵'�B<��4�ݫ1����H�5��B��Y��p�
�a�1�#& �F�Y��,߆Y��)�{f��n�,�E���L�S���}��U.A�Dt8���fE��� �~ϟ��P@d f%?���wdU��V�$mH*��G�,FE^�j�����:�>|�o��w
�3Q0�
o$�yΩ*��o��Vh���5�y��ci��,��,�~�od*@�.���Zz� ��GK��rN�'إ��kI=Ҳ���a���z�~!7>���e�w�n���4�����|��W �I%!:���@u�\������b)���^߫a��$H�?1j����'�~�^h���X��
Y�2�C�7�v������3d�Uk(Ym,�H3��vJ]c#���-�:bQ���nQ^Bm��M����A@kֈ���K��L�3�Ё���HT���׺����c�>�����T�-?Gun��ç����w�V��+�ҒgN)�DT��=Jߋ���~�Txe�ݓj�&O��L�R��w'�df��<x�DyDw�	)b�6'��������g6C�%i� ��MV�=J�cv�$�^���-�yz3K4��jcx���J�[���>�3��NG��*2U��_+ݢQ� 3ZU
kr�6/:�s�?f���4VH���6���:'#�ۏ�^��}Ĉ�J�1�x��;zщ#�w�˥1q� `c������5��[i�i�m+�
,�f�N��#��ڍ��7[o����o��H�?����ދ�A0O�2�ʮnQ�?8�m���Y|f�V
F_Y�Nn��Ī��9|�=	��ר�.�V'��h�5�_67+��t3Z�԰��.���y;�|�5���mn�BZ%�����a6�h��-+y�}�#y<vI
{�XΔR8	`�{"�q"j�K╏O�I�	Gtc�H���G�3���eS 1�*X���h�a�	S.�8���'7lV�i,�pt�X)�3vh�~yq�ê�]}�:�&�03.�5'e=`_~��D���/��Α ǵ�솤C"	x��9;����x��Dw;�D$����K��Q���ً)�i��6���|8��h'�!�ip���e�6�����DtT�W��4����aU��R�
�'i���@/ �����>��.Y^��t�l�S��U) �Ud���C
���6�u+h�w������������6Z"�H"N�	
�X�>�WK5�]�w&N_��65P.��R��O��j�;�N[���	qτp,�AW�n@��lT�4��n�e�.K��멲.6��C�uV��y�s�jw�9�� %���<�6�y;!W(���� U�}|�G��I�31pvJ)#"�f���Հ|��B�=&,{1�.f�.i��a�X���=R@|pm�0���\ù�:N�_�-�q"�Π��&�vK4�*�\�{$��	�TF'#u/e����s#:� ל�;������!@(�.�/qr12�z_ps��B�s���|�)Sz�{fBTkaƾ�P�G:�v�ܑ͆F�!�RF�����k�jS�����I���H�"]�L��~��I�JQg��u�e�N��g�%��A76t�G�"B�-r�a������w8��W����/���-�7��T�t�ln�P�H%]v�$JBM�F
 �$$ֵ�=l���Tt6�.�kR����J@�j+��ݘ�����m�ϯ�7�^�{]�s�kH+X�GJ�)��F�S�'έ�r䷍��%�>��~W� ��B+�a��'�"qX���2<t?DV(�^��f���RiJ�K�lg'�����W]5�Ů����Bzn(a�X1�(T@��	���\�B
�.c���M����ϼӿ��4X���7pl4�"skDb��.�ɖ�L�4�7C#�|�3��7�����{TI��)�(�}����q��\�<���;V�΄qۦO�.�6"�������r �*K�I����(�W�������=Kb��X����i�E�ƹ��������j�j֣�'��r uhZ��������=1dT�,N��Ϝ��4n��ؚ�d¡�5����-%Q�\���èEL��hqsI!����c�w=>���m� �۴6�T�(�õ�5t�Ǜ���(�#O@O��	�Ú�0���D�p/�&j�  �͎�Lus�ϡa�������%HH���\��?�9�S�g�)���<N�\��O���vU&�=��g��"����2G��Z�K93����┗��e���韾*R�H�#��ݹJF�X�G�kr��z��ߢ�߻O��&+�Ê�hI��E��X»W��\a�H��SHsFl��P�j]�7���?�d�uF�hD�B��`*�@�{=I�U�Ғ�L��OD�p^��}�s{�t'��&��#AB�(!M�O���ٮ5}4�/�+�zjO��9���[X�������t%����Q�7/����J�Hl��ؖ?���q����#v�+\	�R�MOݯ��x)��PV��?��F�HR֬�i�>F�s�j1���v��p�ERbR��f�{l�;�p��M��cc-�{��a=�U�.G�\��bfJ��D�_�h�By$��NAO}� �t)���kx�,&� �4>@\V�%�l�=���}��a�=f@Y�D�}�M�Z<�3d ج=��?lS@�� �$D;𗒷���/��l���r*WW>a��,yT�\���������a�:DU6d�A���@(�`��T	��;P��X�X߷�MU�&v#�r D")��:�ءw2W�|h�Y��3C�A�l���F�3X��бb�9Z�kKK�93�Q@G�^�g�s���]hEW�imԂf�b�UzID�:*%�8*fR�?���ԭ�%�
!r�O}��
��)�%��>=L�f���"~�@�fi0�ܺBn���c;��JJ)u.�����a;N�K�<��Z���*�B]����q�� ?�fn�j���&��!D��ڊx��e=#y�:��`Du[�H��'6{*�
����Y�	f�ӓa�a&ƞ�0٦���1C ���7�|���!�jU�V;l�iC��*g�$QT��qю]R��\ aJ��f���/��(�^4�j☚n��E���s����Ns�]��U����@��y+��H��SP��phU�������*=P��p
�.�R���wa�P��@٬��wr�D:X�%
�8�0U��H��Q��T�P��$���[��?���e�%���O� ���&T�X>�_��N�Ce�G��]�sA�g�^*9�Tj�$�#e����/8��nT�%2OB�<=
KO梠��c.�>�y�~��OG�Xk��J�^�s�J���/\�����C{�_D�w�h��7sN� ��1�'�h���g6q<��)����UG�9�d~�KX�Y�i>��Z2;��(���MsF�oF����eԸz��bzH��I�L	���S,���)�����D�6�
� ��֡⥟[��uw�Р�ڿx�}�Y�&�:d�Y�C�����IڎTw�H�R�Mn-�����u�x�Q�\�=;�q���[WWlŁ����:��\�6IW�@�s1#���g�&=X��oʈ؛?�[Du��<%����c��Y�A����p������ ���"�+t��n�"N����'ci#���TXLS���Z�‴��ɓ��g�+z����^�}�K�S�>Ա��cZ�hln����n¤��\u̩�8�Ǐ�Й�+6Ul1�;�v��&�쓖�9x]�e*E�D�;�F�Uym9^�*u#ڳe�EP�	��-ٱ؎����7�%l����y҉��?�\*fG��x���g����O�%����z�ZY���m�M|��x����̳���M'�%�h#����=���s}�-C��
��'��к�q��Jŭ�!�+XPXUмv	�J�@����G���]���H�W圠9���c��(r�ؖ��' ���Lwo�G�Y�5��_�+<�
���ǨO�	�0��'��q��B*�ʚ`I��1�PJ}��.�v�dt{s_���ǋ>�;=a["w"��r�y���
H�OE�2��ț�,Ƨ��Y�;���8�������KN���A|�E1A�N��|��E�C'	�6��+r�����w��,E� l��+�c�b�� Ғ��Ų�\#�̤y��[�{|�^sZ8�{�&����bҜ!�rZ�7Ƀ|��N*<���s��H-�9���2ȨjĕU��3\�]pF����3Y�k@����5g����|�������[�@̉�R�R�}��8(Ú���HZ �wΌ�XJS�ec+���cĤŖb��pv����Υ����D�@�+CC�ލ(�E���9���I+4�,�*]IM��/��o�ٹ�����$|���/}�>[�7�����T<����%~ �bQ8���W�O�"�^W�r�0�wf+���ްT��[�����)�*���*�Pq�9I��hGZ./+V�x�����n}b �Ӓ܏�U�~1�6�f�)�p���?ڊ��$+НY�V~��=I� ��N�w�5�v��O���u�q��wyw"p<I�+\$�@��t������֞N�`�v������f�kR��ic��s�P��Uޮh�p�gL4V����*���Zq����{!J��dG���̆��fTP�����Ͽn�i��Jj�c�H���7�?j�a(��JOJ�p$7	`]�?u5��֥,i4���(*
<�@;�����.�w\\��Kn�~��3Xu{>[�i4�/ȑ¼b:}61 F�"�롺t�l@��K2~z���`z�	����h��S����yg��qH��f�u0"0��z���r�q4;��'ρ��5mq�����ğz��HgU�H�$�5(A�\��Cp��	�5lԦ�cr�J�0�yc���l��ށ�y>.x�V���]$(3*���M~�� 8|bʁ��������7�st��_�k�1��iS������@���seٌ:4�����S��u̡�zѹ�z�D�������l��#��5���gt$y1����2E4��K�����5�_"_~����T�u�D����R��o5���?փ4ˤ�j����%�S^��9p_��q��\ݑ�U+��Q4H�5|}��}�R�"��3{=91r4�Y�.Ȍ z�O�4��^��ɰ3��;T|�����4+`�k"2Ǽ�׼;q���H�	��ܮ�l2�m=G}��z�����z�����=�pr=���������F(q~��s��k���w��f��� 8F���~��H�q�!��o�=�s���c�� /\9�DtC�.L�#�	_�i��~��u'��s$42ƺ�:r(fm�|�6��~[�򎎧��h�w>�tYL��O��L)~�9��oa=�ӆ�;�Vc�2��������(�*�4^����C��L��?���X. �W�	.�	,�%3n���Vg� �x��W,�x�[�w"��*��-u2���=R��U�,��p(Ś���um}.W]>�*e�W�LD�����!����L�H��tw kP����I�G�7�P�~�!t�����L^�x��|�폥��~,��Xfݥ	�K˙s���ztΕV��V�':�����%�p�W��sv!���Q6|�Y��	�����d�[]<���B��v_d��_���>�_@�}�W1e�zݨF�m*?_�lDB�p���g4����7ͮtz�_���r��-��8�nB���>j��XWo$B�1B�ʤn�B�Dr{��yr{�+s˷n5�y|}3d9���z05�Dc�A�i����2 P�(4��S�	�T�ipO�\�Q��L���Fi6_i���!���E�>�W&�H+�eJK"7��o��~������q���X�J���,�z)��^�:A0��P9�v��{��!��ɖ%��ϵV��k���@��ّ(mA���i��_n'�Fk�o��Ȧb��^�� ^��"�CZ�DF(��}�v��@�V!'!�yRdUɤ��d�����;:Y��i�J�+�������8 ���%�Aїmg<���Z��jF ��N����]�>�Z��y�˹�Rv�b_� ��㚖��mw�YYN�� ��e��fu�,�����Z%���7��7"�*�?pKu/��K��f8�_�6'�6ʤ��6����"C���U��v:�Z1�:�w��{%����⪰0<0�+_�OJ�����1bG�-�>�jYC���=b0L�h��^m3��.fs8�p�:,���v�P@.��e���Ð��M�@?��X���dE)Gd[�It�t�*p�-�:#R&b�mP��P���h!��_�:�}��qa�WA�Z �ls�c}]�B���K\͐ X�p!�o��|gMN��P��D۫|���ƆRu���/�Sҷ4����t�F����;w-�%�����y�9�i��uJ�x����	T�C�L"�j�Z0�������%	@�0�e�d}�vafCx'+�9����pD��H��,~_���uy�׿�6d�jl�acm�Dw��䁉<s?c�AB�Bq�Ts��IE���F�W���NA����v�`��`S�T���t�W{��PR�La��b�����$=T�x�G��Rf�m(a�j;��@lLx�'�~����I��M]
��ZH�#l�
��4��X��v����T��ك"��_p���zH���S����"�#I��-S���0�Č���֖'oQ���g��7���N�����_I�{#,;�6��v����W���.N��\K�	��~^k����ٌM'<hEM@VP�K�sl��ϑ����^��ʼ�w�Y�O�s�&Np���ec\��<#@-H�B�`[�r�l4V"��%ɋH�h�|g 4���*&�ePVW��`C�gD�A��pXʶ�j0++��H����A��`ȕHa�A2����e�?}INm��c�!B��K�.����8=w�󍅄+)�5ʜZ�t|�N�Fh?��e?;ƞG\��Ս�$�E�,���_��X(LT9���ClK����VCc늏 {KOpM�V��M��>�?���n�����j��q�-���Ά����54��1�QR����欴��H�̲���e)h����*��8�J0u-�Cߖ�-M§M~�@�I#t�P�L.�|.y���>�G�q�r�Z�͏
�ڭ���;�����qU����^�@ �=���p-g�{��C���}a��<�-L;�=��;�ƁYD��|u')��ة��!#�eg���쩬A��QtpPt������h����ϋ)<Tr�����1�Qv�>�֧C� Ҏ`����o�k�����Pp�ÂzL��5xK��rE\I��r^�N$�X�;$w�����XE����c�I����Fd7��ekdd�X&yO;�ʸS�
Ua�k��(:h�ʫ����1��%qB��>(�O�Q>�I\��ǒ�4��{�F�b�*���~��ɧX�����(�Ec�[��8b������b��.SΣѭ6!A�۱��o:��ޡq�ݶs$m�D�,:@X7b�������ٷy�:Et\Wb؈)�.�Rj=S�Y%m�Q�P!���(EPx���a�0ne�*��G�)������N�Ӈ	+`tQ�'n�&x�{J�S���߂���h@ǄTV��{�5`<�b��x��R��
�X��� kz�}v����!U��Vt��F/x!o���h�f�	ZIi��CI�ّ4��ċ��Ю���Fj��I}\�N�4Y��@"�{�v��2��0WZR0K7��މ!�@)��"m���rx�u�٥nT����PDt��hΕ1ܺ��o��W@Ⱥo=�D*�M�8D�ޡ�szEY�Z���ỆE�R��Ț��(w铊j@�!"I�,`�Y
�ۓ�����i��3��x�s&����|��@q�h�������Q2�$�B��E{��c8Z����)�/�4
���g"Nm� Y�r5�
NDkD�a�}*`�V+�`wn��-�F���Y���U�<�a�J��G�Z%��֣�wG���s�m��VE�ɼ���e瞣=E��)y���y�{12�3G_�f#0��̎�?�IDS��ԠցZ6*P
���xn�1",�'Y�7%LA�
Y$ȽwuC)�@�ݨ{
d?���L$� �bn��}��9�_'�	o�Z��";��{��j�۟w�5c�͸70T���p�<O�f�X�k6Ұ�{?��`y��!���ӯ�t6�.��W��7�JQ/�T��!����uU�������:�r��{�w�,/�f��i�:@����US�A�ת�3���ӓ�[W�Q>٣h���}A�}����>�vZ��_F����
L��r��- A����)��RycZ}ˈ�M����-�����^���_q���>�٤��	e���y/,�&�(�'�i���8)���Į�gu0g4����-,�����pj���5�ƶ��"U�}d��;�p����P�ڔ>RYc�Fx�f����s�P����%���B��݄�z;M���f�w���K�a�\����m�E��m�D�|�j�6N���ɾ�p�]����k�fD�������ա�B��5׌�9o�����ȍ��*f�_����k��I�Q��[�J�#���ٴϵ%_�1�C-�OQܚ�H�y,p&�p-��z��?�rU�mخ�R"�VI�XE!�?|4d�<7���3����{�ÀH�ke��x��}����Q���(n���^��<E��	T9����F��v��q���wP,0X7֣݌��J�Z�%�P�9U��(z�)�6sPqU_
�T��c&�K]f�@������70T�e���E}1����_�& �-����53����{$�Mu���9��
�L[�
.D?;I�	[�r0V�I���	�Zp�uHZ�qգ���U>R<�㺬W?mrGtUB�a�(����m����p\���vn�?���Ŕ6�-&��)3a[����a�ӻ�O�-��kǬ�w��ׇ&��A�z���y��m>;�<�̘`�����+0JJ�V�,�ͱ�
�9������|��"dlz�����������B�6l-�����^O$��|p/K�/(CD�����<�����أ�M>����f��o��0Aѐ�Y�.���>�'q�Ӱ
;d�9\��@��L?X��kAv���,��[�$�¿g�w�����uy`*^����WN��|�M~�w��}�[�p!��im�ǽ$g�h9pfK�9>�^<P���}]|�k4T?t��Aw��&����I���r�ei��m�.s�~:S�~�sb{����Y��5ԛ, 2/-�rO����6�l��1��ܕ��~}��]��Y�s�dkA�~�)��RC,̹^���}M�J����T0�n� �rbBM���i2*r��:H`~�^����UR�Gx"5_.[��m��z�nw���K�;B=B!�BM�G}�hǎW�Cq`2��0>����:�YeQV+0?��[鐕��
���
��31#ߤ�A5W57����k��]���*tR�levd{$~���I��ݯ���W�f����"l�܅��6�d���u���n�M{΢��zQ.¯r��h�O ߋsN�=��k5������(h��
$����,µ��%�����]����� ��i!�B���䊼յ�Nkv-=q�o��1g���v���eߦ��-�05��M���@�5�=�~��jU�;���Ǝ�y�"� �\|��E��b��T��iD��"��c���l�]���{�M�CA�81�n1#���1!�����c���m�,�������;���\�Z`��L��RQ���j���w��gN�'$D+��R �B�b,���(�ҝ��J�0���ln��<>бQڦ�� �(x��S\�轪,0&�Q�)�)���@�(�L�/T��*~��st2�ߩm�H5�/���ό��lp�Q;&��h9+*�'��v�Ҍ"���4������0��8��T�t͕�&ϓ�#�r7�aب��񌂕TC��'{Iy���n�O�T�iLnj�n�_���z��"�zY�e6K/���?�Eז\�o�a�I���խF�sߥ�rqVZ�$L����7! �B`��~�m@{!���Kmm���fo���)�CS������]T̂H(=��c,�XI��v��q��P�� l�V}8+y�C�~H^ ݅�W��n�����`(%��X?s���v0	�=�A�*|��ΰ1�������Ǎ��?���p���i�j
B#/O�`�ׇp����`�P�ֈ%�:����@����bќa�Y�#i��|�£G��0N�n��VP��z"J�dޞ $o ��P2���R7ߖ&(ol!o���6�W�o�%- i�0�nW�c<H��]�AZ�Ov4Iӻ�w!�3�]���
����I Z�9ۨIV��DL�K֘wg���c��T��7!�-S�-7�9���Z��Ã�1�G$�Z��1��*v	mǺ9�|-h���D����;kUn�8�hn�ڣp0�����{ ?c��f��4��&�r�^m��r@���v�V�]H��g!;'cF�`�Ì3І�������I�⥑�L��ZX�����Dܴ�i��)��WaGQ$�״A{��7l�=�ʌy�R��o�����!���%�͆���2Ym%_����&�O�p�Ciر��([5�ځebFg�}l�?��qE�7�a�Z-��<�hJm$j���g�*pD-x7Rk�%���H���[0�$�l��n����h�qagmb��F�ޝ3�D 3��pQ��4�JҾ:��Mm&�$#Oil�ژ:���~�HM99��Z��IM�*�1)�e��;B�������E"N�`����^�	R�^{�5Vf�A����ݷ�YƟ�ij�	��<��z���ҐO[�����ՙj����i��W9r� ��x���˶����Yڪ�d�xT4m�~8��l��H�0Z�;�E;R��U
��WW?R�^2�|7��Eug��� Wȓ�Yګ_�DpUx�%���mp�@�7a>���)A�궶�!qF�%q��A=��T� ��'Ӏ�2�`yV��/����Q-��~��!�D�|�_|�Q�?��J�d�_��~j_�y9�����'�����Aw��.�ǞCi�܂5;�c��ٙ) ��$L�a�7fJ����Ow{�td��k�s�;V!g�AQ� Ȕx7�cU���	4/�f�]pA�2���w+~�!���#I'���>}�Y�ɻ���:���R��>���$��;cY��:�O�9��΃�sP��N9�@8{/_�L�R���wO�ni4�8�R���c�4�M+M�6�=|r�е�%톴��u�u�5��r�t�8�f�wIH\8��=�L7~Џ����@l�cN�'��W�c���CY��d(�`]�N��{&�&=��貿!2H�JD�K������?)aM*JR4���ӹh�䑯zsSp'�wJ��noR�[?�|H��� �#����XF����oYxc��.��`[�~�x����O]a�!��zt����DYސ��y��	2��]#���	Z�x��"�K��c���,ߦ!|�d�bt�!�Ӥ�������O�ٽ9�z�\~�-6��+��ӫ�P�>e���vS��P(X�j20/b��m#v1����<���q4�{(��K�"�n�@�t���&�"��Xp4��a�<$��L�~sΎw�s.��;�N�^:��j2�YP����g*�`y2B �10h�_ȣ����������=KzxcM��]�<%y_��_0\��}�5��g��9��>7���<�t9Z������+�ơ��q���p�@Z�ᖃ����FR5���q�*�f�)1Pnn��
_��z���1ynu��2��=��yQ�Lej�1��$|z��P=]ȃ�ΚS�	�ȹ�jب@��<b pi'�����z|�з����t�^���D�����U	�27��EF��F������2[P��hқ`ˏ���b��X\��J���[�l{�P����J���S�_޵��2 �B�6�j>%���Ha��X����y�@�f�������k�iP1�����Mbޕ����RBe���nx��\a��V�և�1���X��Ŭ�����?���'ĨF.�3k��y�G����I��Q���m��Ë%�=����snr��BQ�Y��P1��&�F����-"Z�0��2��%��t%�(��.6M�� 6��h��}H��:�̏�����ma��a���-׊-�)s4P2}���MƳ����Q�T������	�V�	D�M�#�iW�ʃi�������@/0JW�{���O<0���O=�q���"��;.ʁ OZ��Z�n��Z2���M'| Dǲ�-�_�'��@�=)9��q
���#���_2�q��K��g5�f?c�Ÿ)�o�7��\
 �������{�)�3P��q�W�}F�Î�t�i���K��w��=6҃IpP~.��ғ{(�I�\����{ϡ��nw��8{�A4{��?�@f�gk���*կD�?_��m�2�\���#���[�_�E����Ț���͌1�דϡ�"p��jJ�0��yىP�-ɓ:~y��{8�,��r�F��:��7Д������T]��T��#��FU���H����<�(����وZ|��L�3��=E�n���E�-�ᯡ_���񚴥M��|�~i%(�r�eo��(.`G�1w����#,9� ����K�Ir>�z� ���1�]���|�i�����nJ��yN
m�7���^�/K�+r��UFZ	:�Ҡ�-���.1ֆR��/+�^=l;Ҝh�j���8�)���4Y�{!C�
��Y6Bv��������ܼ��A�s�5�d�Oa*��GaV�T��#�l���p>eCNք�Ҳ��]�~r7�(�VU����2~N�)�x���$.4yof�g��Gǃ�Tjj��.Λ9�~���5�GX�Py��V��xA��%�������_��H5n�ݵo�xzQ�ڈ��˾>vQ� �M�����rD��⢨������(*Ԗ[�PZ��<GK�7��{$�.��Y$�r���,I��_F�;����N�_����٭��^>�>P�sLʏ\�����׾j6?I;���X�`9؂�7X�u[��<u�`�ڨHB�e��@h��̌�������9��l�ذ��1�N�Y:��p�>�t�Aa��b�*;�ð/Ғ��~8�q���!�s8�wo��c��3��q'�/��a��%'n��3��6HK �S��\�e�<�퐂��c��_�ү6�H�k��v��H�L3ܔ,��"��S��dN��
&�"�1�!1��]_6�� .����Rr0Q��~Bӷ�1�_)�{�Ol��8p�Fsn8�	~��ծ� ���,ܕI�+4 �#��'�	$��w��5���@z��.�c6:�mu��@T�������� ��K]Or��=ƗK��X'�23L�B3-j��X�l�	�G�]!����ys���x���v4db�D�~Wzg�D���|�Α�2�.׸?֓�z��x�Ylж���~��T�T P�Eө��_���c{ߋs��-�b�]DN�D\r�Żn�س��W7~�:�7��Z6N�w��-�{&W���B�'�+���f�qwةܞ��8kT7���a�eI�̙߬TT9�;��I�*�pꝐi��	l.�J�ς��9,���_�3�W_T�#)�oQ�O��$kx�1�͢I�k��M���x�0d?��2Qi�&Ll�t=�9��64�ɟ�-[�{w;e����5� q�7js�����M���
���a��ПC�`�4�g*�J�y��r�M��{�zuq�[!w��� �j����r����ߡl���d0�� ���5��A�.������nbEBw���YH���@	3`�*����~�z�h%�`�5{�=Z%�ͣ��f�.�7�LZv��_�Q���d��1�Ə��E�λ+�Xt�̤
V�d�I+i 6�����}%�-��$>֕Ma�+t��_��+(��̎�P�D��Aw{p���n\�9�`#d�k�V�(C�1�^v�m�T9vw
�؞�;D[eUZ���Ml	8X2��@�<�g�[,Eޱ@e��%���$V�b�,�s^Px�� UJt��D�衶x�=���<�1=P(�A�窪Y~�hP��)��n�,�����c_���n"ɫ�jȆW�y�H?���e��_Z�}�j�z��O�Xf1��x�޳��b���ץ�.��õ篰F�d!9�E�߳cIb��3��3�^�)�Aj��:W��#R�!�:e��K֣T���%�6��V�D���:BS- \F-k]'���i��N6����0����G�<�j�!��� 9� ��$S�_~���b��U��.�:�E|f��YyϤ��2�c���:��T��2�s���宊bF%�G���R:�JO�E�2��uج��O�`����V*���k�K�E?�]�0�޼&8l��m���Bⶵ:O7�`q �_I_��16�9U;�#D��F���t�׵��&��n0�OH'�2�]I�����(v��¾�C%˜~e�@Bww?�V�W .�f��<	U!��ex׮D5���`XL2_�tJI.��`q� ��y��ԅդ����H�&-�&��wg;eU��h�5Mw&�n�K��g�3���*�wy}ӗ�A�P��>>n=f%�!���,Ⰾ)2�>�'�,�`+���A#5ޏM>�i��Gp�>�ܖ�Ӯ��i���(�.��T�!�7W�)=^qdjf_����� �ۻ挊A��J�9QV�����80Far�M��4P��څ���(�P����F�l�b�$w�{��؉�Q�����2�}ɱe=����� �2�cf���b3KV��u΁W�mO�@T_s�z��m\W�aD�U�!�q�����t`��i�{��膻��R�����+�B�~��3����r Ȑ]PB�����|(Έ��K�u�F߫��>tu�MT���cx�
�!�'o�ټ� g݇�8���`�B#s�>�,��ʢ#l�F�L��gA~	�*B8IFLb;�O�_2+L@q���[�@�ɝ�}���.ԟ�2>9ܣ&���o���6�ŉ{#V�)5!'P���;k�C\(	��흆���+?�Se�Ø�����E��C�UAB�^E��EG��t�M&���K�M�_,�c�; >hs� V�r�h>��I��]pț��"'���菁	�B�@���]>��췅�.!�a*R���i��ρ�@��-O������Vji0��h�&e8;�S�ۼ��cnZ�a���0�2�(4t��Y<*����uy\�[� �5��9!��p��$��z�t�@u�sS`�IP;Y��ƀ�:=��s12���6?����{i5�$����D'>mAm�����l����qV%�� �"��jg���H��6SE5���X�]s�5#��;䆘���V�[u�6=$���i2��K��䩲̎C$�S��RZV���jE>���ax�\�K�A3x.ĸۗ���U��B	�I�onھfgC��ϰ+B����t��L���P�mQ��2;O�rl]��e��S�K��ݰ����[at����:-���͑3Z��Z��6��N�{y�� ���A�m�f?�� �/�^Έ-)��Dy'X^R3t�X[Il[dg�|�/��o���8�Ij�9˅�a�d�6�'�$��&�{�%7�%�����TF��TH�
�h�1�!�#�7����=C���2�M��m�J����eT�͊�L3uyNO���B[��W��lv���ѹBKv&Ļ�H�
�K4��G'�V`��Dm�=�	�O�\����u[�Vx�7���nє�R�'bE:��`�z�p�w+;}��=�������D؇��� Z��9����7Y��ӿ�VO!3�Y� �'�>3��BW|Wc�;(��0�@�����_١i��2��X�����W/��
���KV_~��\.q���!D���G���)dH�'dk.um����;n8;b�w���
'H!�M�����c��-�fl�U�S�G�h\��<��"�gZ����Pl$f�Cd��q���^�@@e�g�JOϩ������d(V䓅~W>��C����%C�L�?P+Ķ���<����{��ߍ<
1r.�2(/B�{�x�T�WJ���^ZB@��������3�4��FDv����y�|��v�u}�N�q��* [l�9���7k���^������nJc��>��;��=�R�ɥ=GjZƀ�u2k��r��Qv��>���g��>�H��k�lKa�@��][��˹)�~� ��'�#rK����XwDД��tb4�a��(�3A
���g�.D����-���D>����g^�PL]�]��;��j	}å�'.�8� �b����8cn��k�<;�O��l�F��I�w�p�Y8�q:��̱�\���]�$ۡh��<0^W	6��̳_,*�@���z��P���&�靓l�|�^��9(�2;LɂEi�IP�S����[���U3�į槫w	��Ja���2�fS%3��E+���Rb��Ԁ���J�I��F��N�m�fZ]�7�Q��eV��m"̾<Ab��n�J,#�ÌJ0�1��P�/�[��Q�Z���/E��'�IA�[J�@3�W��DEB�f��̬c�ڴrΞ�YgQGŏ���Z�7l}�]*>��H
��ewˊ�
g\j8$��K��7b�fAz-��s�=�?����qi T�F�/�$�$
�ax"��G3̬�j ��h�����[zKpD{ܻKMG]8��Z����������������7u��c�����6A���g�m�\6�� a<��9���z�s�Ӹ�;\>s5Kr�����C\$��~ŕ���� ��!�CΕ0T���uu�ER�.'���_ �nn��J�r"���ԛY�j�g���h5k�Ԋ,%6���������,������3��G"h��T�+?VOt?��
d&�)E������n�ڎ;n�3A�\���-�d�^&���*�yl�X�{
����VJE����q��)��ϕ�x"���`��xY@��4�i�|��E�8bC���ޟ�b3W�,�� �JF���F��g	R^Yߠ���˦a�d3�M�+�H�!���&�:2�a���.�%�=}���/�_�^�٭��Ȍ1��p1��X�ߟ�i�2h��Z���5��$�r	�܇Vg������K�R��>�-�
7����C6����8�B�����5Z���J±�_�2�K)Cֻvwe�h,�_Ft~AF�.������/���Z�S'�c�X�F%�-u�X�N"`�Q@ބ�Ї4dD��]�?R��t�� �*�}�;--�K&a�y��� �R k���(��^L2=�*� i��iCRA�	���9R�CMܨr3*7r w����nyp�&�mLx#vl�%갘#�3zyg58B�!f^�'���SͻxD���VY �[L ���F�;8GȐԪ�e�4d���޶��p-������PA� j�^��!e˧-�W�EY�3u�-�Xw��Tx<t7; i�z�y��A�D�;�Z�Aј(�j�	��C�O5~B�զr>=��c��s�� �U !�ZQ_h�I8�W*�К1�E<�L�۔��>��c�D�3#O��Te���K�Lji֔TJ{��*�r&5.'�B�e��k�����^�W��0�M�W	�	����1w��� {��={��"v���tS1�����!nv}E��*?��x8b��d��-t��q�%B1m��Ϯ�N�����sl�?{&>h]s��v5�<u%���)_.�'J��d�,?�
j�-���#@00!x|>�|&c"rx���Se�a��q)���êh��I�2lie���!UI1$���D��@z�
UzgW�Aʰ3���OG%y�v��,#��:_A��$�?J� 5�MR(8�a��6m�iYe��Dxe1�~�I��!+��O�]Gd�56��g��BXA/X8��1x�3�0/ٍ�W��V##o����?���za^��OƦ�X�s�O�~o��н��v�a�ST�h�|w����"����@KI%Bp���K>�F|�&6�,|��	8�;�J��e.E Df�C��kCY��b@���k�Iw㻄ӏ/�d0 �9=����rq��/�#>�rD�
�|P3��b q��)�M�(*"��	�����3@�VW\]p
R�ȅ����B��:��[ �4�r=�4��S��:Z���v7w��,	srE�k�j���
C����+��A��L�OSE9���j<��{����uf���*�@��Q��ÖX����~�fHչ+��l��ͬ��š�HL�� �X��h�o���:]4�1����s
jqUMw
�r�'����!�/�@;&��t�.�kH�S@n^xn��~6����6����D�P�VH���E�����+n3�7`h �ƅ�JRL�dH=��yu�XG��+�{F�zgW��z������/b#�6��,����G���� 1�$���}�
����>AYŐ�fT�G�e�~��]�!��5AU8ܯn����j/��хW�q&�1c�ȟUs!�+8�t�xAZ^����Sz��5<���6Dx�t��d耓Ew��i}6y}W���~Y�X<�oa F��"*xN9�dA�X���7�np �}���@8_vA�FJ�	����w��P_6���G�,���m�6�w��WǶ�����>�"��x��	�V3e�z�;W���,��1�3�(��eb���IE1�	w��Z�-1�
h�uٟ��>11Ү_�6$#���D�@!Io���2�Rʅ�BJ��RO��g'X-�A�'Im�i�͋p�`��|.w�i�b$.��`�͵'��!��������=��*fr L����C��߇�϶��ү�Ӽ���u+�ֳ��p�dL��G�lg�Cg������t;l׽��~$9zD�;����O�T�������f��2o����`�y�D胎v�G@^3����d>�N�X��W� 1M�17��HhW#�0m܆	�� ��%�닭�-ӛ���\s��O��[���Q��~&�9�9���Ž�iK<~���㪿P2싅��7�F'J+�gЙ���`[a��-�5?)��z3+�V�l�T�P\E��;�'d':.O���V�*�j�`��	[�R���v�J��?e4Ny�=TS}�d�����"�Kg�������
%]��?�_w�I	��׵�B�!���P4����ꖝ�?�v����$s[ƣJF�M.<_vE��-`���V�N�>��W��+�[���&���bP"�W�kC\��K�1�0c
�e�JW�[;(sj �a��\�5Y]�]�=���f��ͶJ1��\�k�����TЭ]2��-He,��÷ك����S����<�|ʃ�^-:�;�N���i�ϣ�G@+�T�bJlÔ���?v�����Ou�M�@���K󈓊&��'����s�i�e`(��%MqZs��$���uK��$�������k[8�����������1#��)���{JF�:�������W�/��"�u�Z?c�����_'���ⅎ��[�u�U=���o�?�
B{D*��!����`²�.Z�w8i��$S���H"z����������%ɥ�_^yH�2��񒘕q�"���D���D�=Kȯ��u�i�W/�Nnr�bq����HM�83hU��IV��W)�F,g�r_<K��I�ڮ��,;�:�V��]��"�nj$2���6��3kM�%1�8�9ݮ�g	Qܝ]0m����X���9XLj8� 3�vPC���E%�A.��e�^�]q��.��/|�>�X>͗*��y��=	$YS�jR!	�@@>���~��\���F�����O�N+?�b����N{d"0K��ш���i�M:�����s ����C'|���@�J���o�c;����p8\��d=�2���}+O��Y��(nY�;�-[��u���c���b�ߝ�F�巜K1"DMj�Ll%E7ku���нt]�o��Hj�[�F ����k縶���I�zv,��@����\�4p�#�q�䗘�Qĭ+�'��PP�t�'Q����n!�:Y<~v.�ʃu����[�o^�'~��x��: ёd��:�T��A�E�*�GwÉ�b��^�:���$V�X�/u��\���8�P5-SgP>���j=�sI��!$�Dz؟n�d-�g��-o���U"��674	+�].�"S��fxM��%H��}��Δ�w��UF�>��^�:���(�3YZ����/����My(�o��Vw��	ؔqd�%�q��h� �m ���FF����<�H4V�ao|w�۷��fVH<����J�l_#z� j��*LaO�T�� �C�|��ii�2A���B�}dX#�����hp�H�X~q9�^ޥsD�Id	�?]�����7?$D�0����9N�F�d��[�M���	�����"%���V!��:�>�� ʾ/!�S9-]~��i�D����ZÞ)9vFSڷ�ݞ7��g<�?�3�vN��+~���=���u�,
\��	��	�Qή��32���Y-���픽�T֞�Kn/ ����|�'x5��x>ԅn}גr~3r�;}�u̸a޳]��yCfl���a|K�F=�ϲ��Mk�m`З��n���2��Ɏ�72�e��\�̸�z��c�4W�u&B�w2푡�H֬r] �C�0���t��G�t���ۤ��/ھ���R�Btѳ�2;�-�M@ ۬S{vf��E�R�:�"��p�#��[�M��8C=J�M��"l2�W�G�7e���W�9>�J��r�l������B�`���h�:zpL�F���5e�f;)��Ҥ��̪�t��!�1UӠ!���riY�WL�W���b^�M���į�ɛ��iy���F��aW�H�=M3]_R���[�!�B�\^12��X��PL!*(�.v��q!��Zc�q�� %$we�(��dY��Rt,�º(�e����xp�_nt��4�<l����g]���O����n��K���Ց�/|��J�8������b�C�iFߠ���q蘷���ݮ2?g�7����M�K��Ý�.�]�l֓�3�H7I��2W���Ȕ�L;����d�{��B�c[ ���S�����!�hscRD�>�ƌq֝�V<�2{^��#wn.c83p-��)�g�fC'ֲ�S�A6�oeε���y�eJw���#Ҋf�Ta�9���0�A��'{�y�YX��	v�q�O�i�s�Z��O2��!}ͥP�	ۧZ�6��t9����V��7�}�o�Ib��N
&4�ǖ�M�/>M�xq�<o�l�z���-����:��BK;Q�a�����_C��~�F�)[v�,�!;�F��5��-O-@P�6��˖94����������%�ԉ��n��O��z�y�P�fpow)
n�̇I��O��k!w�Jv�ǻ��ОgZZ���;2~݃UJ�>_5W؄�_x������ն���h��4���M �n�P����M��X�d���Z9���n�<�ȫ�ȍc���Ɏ�+<�ں�N� ��檜 �rX�j�`|1��KF8o?E��r��	��~ք�s���˳ջJ�i~�@�A!��吟p���qo8�.v�a���S�Q�Ok�{�Z"���X�&��E6q%�<��̒RiaU�@Ơ羴��ݾ]�/<�T�j���գs{�����p�|"��>os}�>�D��;)g|L]��b�S�-O%?�Rǉ'ώ�75�S��/7Ĵ�7K����=w+���aR\'�E|!&�
�Rn4��;uS�����lA5G�a�pG;%Z?C^�C�Zb��)�^���S�n��E��=z������_��SC���-��()�1��*V/j��R<�@�� b�DY���{q-+w1��b�!k<�S���J��#��7��&h���]&����[��-8Ʒ\�A*������<�M�A����@�""V\����QiKH�$���[#5/�I�PՔ`3)L�m�	�� 8+�օ\��C�I�p5c�����_�%�*'M���������껡>?c�S�j<���9�
�&��K[8T���g��q�p��RS�Q֙�� |���Y	7�+���㞅5�@p�_St~B��Flv%AMuV{M�egl�m������	S9��8��T�����l�B)��9س���^o��w�#��s�|�gD!���|te�����t4�%4iJ���%8,�wy�I���g]�lZ\���;��G�08��6��}��xknC�e<�X\�-����K��: E����S*$�Bz�S&Z�Z���2w^��M� x����g�0n�st�H��E�M���sT
�d޶����U��\��|�wM>�0����X 
���11t��S�=�]Ha]����rU�pSL%.�9�T,����xp���-��^�>R��q�uy�����{L���k��$�pL���m���3
~���:+�#��[��ۖGm#�w�_�T��	ʚ�6�\.;/	G���3��Zƺ�v%��o��בy�UL(�a���ۦ$+��$2~O/�6'�*H[�>4���(q�9�khGު{�H\~ut�f|m�d�|�
�qH��v�\"�q�f�w�Aуn>]W`�����*�[t�0\�>��m>L�:fC34:�-�z2|y�;�d��x���'���<��?ߕ��nnA�F����%��M�E%:��Y����ێC�#� K��r���,��N/:��R��:�GB��Vop���<��L�6*�����\J�u�|���ʙ�렂Wk�5�m�_��:�5ޯ:V���w�:%51�>}���qN)l��&�s��k�x�0�0;	T�	+��T*�`�@�CL'�� �����ƴE��@c���ʶ�-A'�[��I�Ur����G"ODY��f�H��w$� Ɠ_۠����A��>Y��f0��܎e��Dp�D�J�K�S������1���	��E�&����R"BA���{n	:�^3�N4�3vO�/(� ���5��c��E����ō�/�D��d_/�U0�����tʘ�Q�{��.Q⚰�����y����,���p狡���Bl'�l�nVQ9���Ʃ�}�U�T��������y�1G�j�8�P&���	נ�WMƦ���L�T��SbR�Ⴢ�V�&#�$����G*8�����x{~� +�FWr�ė�O�a��5�����C�3���J�U6	��g1(�P�<�HDkH�� �5t�XP��a]�_�V���Z х2?�B8�e5y�+��R��o�T��0fe�bK�F��ߡ%����ț�H 4�&Q͝��nrl��[^�ǆ7dǠ�፰��'()rW_R\+���C�H�>\�|BJy�5�T�8f�ֶ�6�Q�YZ�X,�8���ܣ]�d����k#q�'�r���1�z�P�Q�~*��=�'��Ә�����8���+�گ�]�VG��;L�u=�O S�m8�WV���l�}s쓣��� <�mTmM���~
��M����{� R�䗱"���d)�����<Pz�!�*�&���3�Q��%��q�et�9�1�^�Cw0�;1v*��\f�;���Q�IH��i�-������Nl�(�(=���
�v��OZ�$&�H<`Xn�f�.��+@j����i#�5�LoG�@�#sF�l��V((���n�� Z�5��f8���I@�DvD���et�}F_{C�=om�2G~6$��uk:�V=��tQi�N�.���<��O���D�I�Vհ2�y�UC�b�ρ4��m�M�m|�T�d�p<���_7�M/�L������-��eZZ �(��5���@��]�p�mc�I�\�]�xDT���X��_(P,R�X������d�C��!1��A�\Qs���Bɢ�P^ ����c3����2�>F(��m��P>�.[2�K�V@�V�l�T�$K�9��Q���ϝ�|w�Bi�`)7˧�0�3'`R�4���%=���T0դ[��Q�3b�'�)u�͒��O�
�q�s��t+-��@�����������ͤ���k��mD�Y��\`��NssL�/Su_���,]��^6g���gOA/��1Ec9�����9;�uy���˧v	{4����gq����1O�8�;����{aY_�f�����k�	��E���o���:p��i� w*�&lr�XiGѼ�v�P%Bi�����yE};�O=�f�R ��:���	QP��*pݱz�4ƫ�/Q�H>/�E� Err�Qe���@�����y��j�ݠ�Xs@q0��a';8���Z�t���@�R��C:�c��~�2���*�f��h�Dr9Q⏅K�o9q��Vs�S�d�Kn���z����y��ҎQ:��d/g£���M��-d?��+��dVH6(�{�I��U>ݷ/�#�1D.��Hk��rM%���\�
Y�L�c҆�>����oV����w��)!X(G�r� 2v��1��tNk��rG}��{n��<]�����
C�2��X#�C��B�S:{uR �I�����H�ˠ��cՑ칺N:n`^tT7����:lS�_�A���`\���誾(���dۖ�r�٬�28��ް �V�����_)�Po"��C?&'����!T��h[�c���]RL�:y��o��g�Ώ6q��N-F�ԝ�J�@#52�K��d�ܼ��z�f+��c6�������z�C	y�ip/j��(�eF��	4���!��#؋~6F��B�ʹ��<_ه�Q�؜��A.�Q�@���V�xU���~eZ���u�D�iz7U���d�� �P��2ʔ����Sb]��ßz1���)o.����b�1��+��p^�f~'Q�����(�g��,kcmx��9�%�;#��j]�qꑁ����.U��CM�UE_����_^>��ͺ�,��ƾ��6 f�cQ�DqY���6�$Ց$XbtC�d�n'�"�����N�{^n?�P�z�����t`(��T��q���y0����_��w3m�7�;���"�4X�Լ`WH��N}����6������d�c�8ш�=$����"=z�K �0))p���2�W6%j�\����a$ĖNS�{��rѵ�Y`��HL{��=lwE���vw\P����Y���c����8���@�P��%��w�	w�̈:��ҿ�:��h���-���̸<�%K�a� O�qTf�i�6t)0��<�>���w?�
�$ЬO�'!3�`�*�ͅ�Ow�\8ih������V�s�	�3e��5�^��N
�58���Ro���*��cƍ<z8v��P��-.��S-M`�A!8�Ȯ�|ᶄ@-H2�!�>����_�Au������V1S"�0�e���O:�)m��;,V��/ZM(Ʃ���0n�8��2�Pn�� �Sr5�Y�n����N��hơg�U��k�Ajs�*kW$@t+"8��4;�9N�R�7R�do�Ŝ4'���ճ�I��%/�Q���j��?��nE+9�uC)��iZ�^�S�t���(L��
���T�0H�#"����A��l����}�/yI i�ғ������o��_�%���F����(�2�W�K��
`�Dt�|��T���C�(La�z�e��@˓Bo���c7�;�
�AQ��V�o�m�V�z��B$��SGds�}��13� ��ߎ���V�s�+���k�i!�K�>.��P�%�ٽ�dm!j��*�Fd��*q���?,�j��}�;��<���st���A���`
�ħ*庭&�i�!�������pE$U��p�����m(�Q="B(����Z�dn����*K*%�]uvV��^#�]b�m�aX�2�{�$��D��_�i�~%�U̐=�����$D��Bl1�v�U��}������}�Y)+�/ң�./�>�%E�C��*�KZ��
���f�dhw�֬���i0�����uz�M�P+��rm���R��M��V��MY����\��̙���>���vV�r6aǱ�Ì
���'R2A��
�b�	s�޻(V
te0}����&��N}ɂ�a��F�wiiغ�]x�z���Z�<�����`׬!εS�N����-{�w�?rB�3F�@���[�3��5�\�`iyn�9�e��{O��I�1�%��W���(r�՚���:	����@0�T��h��D�w��e�v�:갓��{�Ȼ���$�pl�#m�I|�Zs��=l�l���0�87���tCj_����(�.+/Ɇl�] ����;��Fbq����f��b0�_��
1�i�8sj�*Y����l'����̂50!<���N7S]��f�7�.N{n��[�-�um�]�H�1BdDe;Μ�3K�o�����EP���C&Ȅ�u�2�ϝ?ph��E���j�;ݣ�#K�g��ݺS,�@<�����^�,�5[#sl����G9_K�8Kn�n`�[R����`�y潻�FIPmf�S�o/��x�4�{�&u�Y�~���z3��5qIz�b�e	�(��V�f)�$��ۼ�m�� �
f�y�EV������d�Q>ɋS��� �;�;��Zt��G&��¢!
���G�}5,��D
���r�R*�Id��5
�o���M�4H�çIe�D!��3HA` r#�}��q���0��)��VI��Vq����S9󑔨,���b��=)'�# ����[~:�WN-X���j��@�V����΋<�*֣�� ɉ�V�z���� m�8
�CG�C���Dwq��.�Ch[�ޡ��6�,[uDBFQ)꧷�.�|����C����Nb 5�Ƙ�'�Edf� ������C���ɕ ��F*��*�L�� Yk�Fa�������ju��D:C���`��"����F)��<s~���P3�-~�m�v`�&`�Ĵ�o�a����la��0T�V��Ϗ�d�Y�G�`v�bxj��m���`���:� 9�Fz@Z�!C��yzp7�G�7��z%��#��6h	k�]3�6ܪ�`�I�@O��`w��t����u�'���N��I���i��jZGl�u�<��MO�"_7�M	,��Y��F�"kBj��F�v�(�o��r�7-���g7��L�R,�'��2��)�~��*hU&��c	�u�$δP.(��+l��R�:7t���^� ��O[�ޯeP���l�p��0��#V|E�XY�c_9��̌O9�C�l�w12`�����Y���+>���x� {j�6����l+�p K��IA��S�
6g��<����3��RKH{��v=��U�:�>�Gӯ���$�p��۳7��X�`}�o���"�����R'�8�l�#�}�}�0	Άq
ӂ�#쳬Ϛ��8Q�kQEГ�1r���EZ���]{8%����FT��ődfd�-6>O�"vxusa(��>k1�TK��8j9��ib�m�L��F����{>���*�i���˻K[�5�"��L�N�R���]"\H�ԭť��?a�D�_H&�r�
cH���?㛥�r��{k8	�/H�%�)����������{4���M�C�͹0��W���I�s-��^H~�����0�J�Ur��$���1�+^�++��/�ܧS�(����,�o��7�� ��3��֮FL�n�̕N@D��4��H%o�Um�����/���=��ȋoZr�`@�'L�����$���;�����*1������yfN[og��p;H�o�I1F��Q�j�!�յ]�[]��}z*���M��1�A�K[��)/%�W���R ���_/��Yb����#6x�P,e��9�ס"�%��W��ʘ�j��,���v�+�X~���}����e5����k��>|�yT1���͗mdo� �Z�W9���4f@���B�-�v6%G��Y�ㆼL.}��f���>{I�J�ٌ����7@�8���9yn >�Z̶l_��af����+$ ���T1Z�Ҁ�W�Q�cRӸ���
��_�Ǻs�8"Xzͱ1'2?pG2��%x�R��Q�A1���o��E#=��ީ)��)�,ڃֶY$NI8}x�XF}NB��^�E!��Y���*��(���{���w��В��їl��	��s幢��?�1�͈E��@�2;�Y��Gu8<��(L��[{�?J�Ӵ=��'i�:J�ʮL!�4����:�4�E4�,���q+Mܴ;�FC�Sz֑�W��+Q9��΅i��0N�����Gu��M�گ�tS
�-Fۛ��9+��Rj���r\bV{�~�$�@�lpzF�J�6�y�L�|Q���R����
흷�K���o�/��r%M�j�1��,iY��"�ZW�Y��j1�|��f�e��-E�֊��҃pAޢ́H�-
�_���3/z��+�(=+!�oD�R�_�р��o�����J�z�Ue�dx��V6����g᭔]"0/&�ʗ�Տ)v��V=.�5n�4kQ�o�KүO�sQ_��T�@z�B�X�C)�_P$]��+��|����L��d:��L��8�>��T ��N�z�<�kqt�l��9�*�o���x��T5�O�u�+0���J:�m�`�$��q��/\��-��gi3�9澂�p���Ab�y>�r���.�A@z"R$�詭��D�?$�њ��Jv��>m����.}�G?��~������Q_�5�i�Bdk��	�� f'g��c�4�n�>�����A���L#Wo�Qc3F��u	>0��O)�:7*k?��${�ׅS�7r|�Z�d��@�����}�;�|��%���4�)���od�$��k�M
����ug���>b�N۲��'�M��v���*x)��ְ;�w�᳊=�]'�8��%'#��<��D���r[�V|�TLvP��ײ����}�V^!�=D�Cy�yG�.m� U0���h�e�E��<�R|��r���+�ϚK��`;�֙ �G�h���jE!��_����!��s���,�7�ͩuj�`�{� 
��KHbG,r\����K@�)�=]6��� ��F��.�N�R�DGJ%]O"��Uw�VH���#�r'�T�屰:�����$ę9�V6����/���h�IX2���[��i��X}Nes�=S������mx�ڭ'�$ٵ�g��e�q��|C��rV'>��3"d8��k�O�?2ʗ��Wb��/�P-ы�H.㌞�|�"�ɂv�2Ē�N�d��%���S��z ���W�!	kr[{*w{��Q�*�����v��g1K�s����[�jmU�9�t���9o�� ���K�ϩ�����9�\�@H���w��ux,)ic�'���G�.���t�χ���v �o��m���,Rq�l7���%�}i,	6��(E���������3��v���[g���8��|�h�mh'p2W�(�(a�GS�s+p��5�b����.�����¾��V�t�`�����W��^=��	_HXYݚ�#AR`���gI���,��~�[�0�([3�yvs���Zq?�&m�퓵0w?bu�,b�}^E!=�D=g|��Y��҈��ތ>bo6=��-��߄T��[�;�28����xH#נ����p^F}kL3�g�.Cg��(��i]����b/��nQHap��^������%,猰��b*�!����Ô"n п)�Z�����:�u?+�� ��=Ls�j���!�w�F�3���������hnMU�ª��G���e6�te�P�^j����C����:[PL�Ə�N�wטPi���5��m}O��&��Z�\4��vt�2Hc����Y�� ��E��v���%�fF�gu�.�a��DB.�e1&�З
������'k���r�P�ˀ͓�U#ɧl�
v�uz���Ǌ Z?ú�G|��gN��Y������-��"^��n��|ƑWV����I����G���y��.t>�;g�8e?8���vؚ��5�^�(�m�S} �
�F1Q6���1�*x�HZ\'͈$s0�fA2��m�h�\�_���O�Ԁh�$�?nx������4���8,&>m�-zd�v�� W%f5�tHFMo,a���i�CJK���	��%���4�G���#k|�3���� ���Θ�_�K�{�I�� A�X_{�IG��[�����#�:A��d�]@*�?���z�Lq8�`~5�o�~�9�y�8�Z���M��ҿ9�!�2��x��+�S}|I���V	�m�릀)�&ta^Q3�S,�Q&��I��x��]��5_��� �58���gB��ͮ;rY��C����5����o0έ����ӊƆl���U1��޸t'�{|�j�:�6V�ONɗ����y�A8{���T��g�+D�c6��I<�V�+�s���F�@N:��fzeU���ҥ+7,������?P�uj׶�謖'�L*E�'�hR�#� 
�<a`�લ��BxI��'��r �K�V���<k��eĆ<2��7��l7d��L6�,���7%��8����>����#�g�^+���s5J����c����8o��O{������8)�����c�lF@�e��IjZ�D��4H�E ��V���瓫B��ˉ��í���x��5���}V?������'��f5؋�<v`A��|�O������s~����u�nj-������ߟ�P����/��o���8~L\R���\ŨV����<{�?f�����V�O�SXD�1�`zY���&L~?���k��F�יWV+�9,<��t���f��pj�<��3\S�(�'�G�����6�5]��'�c����'d<�q��z�O�l���͕�NΝS���UB.�|u�ͷ� ��d)bsBC`��b��.���R�WB����2d�Dt��bF�C=�'�?�94ڒ�@��v$�J|^�,��Oe~� ��ML=	���F��Y��^c���Z_��90i'�����U$�>7im���'g��q�Y�)=���{o��h��H7��Z��f���������&+4$k��fX�}m}i�����H��7����W�@~d��GƩW�J�0�)��S�WT����
"����	����.��QN˰V?����X:�;�1�V5;�[<SF9���`J��ơ'��.�T��gLF�	Hu��^M���Eō�)o}\�J(�{�A���d)KՂ�Ӎ���(n�hH�	��)�} �O���V����$%�N���; o�M�����%��!��눙��M��Ū�?�P���]�� �ꚱ�܈���A�נ4hs��`f��˔=��~#�hr�1��m�!^+x���0�h��$Ec�J��"k}e*O'ʧ�@�9�9C������b9���}��e*�K���X'zrg�}*�-]=�/r<�p���,nk��<��a�=2u&<-� ������_�ȁ��?fd�[Z�ڗ�����9�[x?�n�n�ik�г:�TIN��N�u=������ @��Jq�U�yUj�c�s�%N~�KZh^ӭ��bȣ���:�	�����*��B�<�֤)D�� %Aѵ��+���fd��~�Զ���V�� n����H��3Cv�08nx&S��ӷ�F����DFPn%o�yH3�)'����;H���+����J�<V���?��a��DΕIB╣�ֵ�O/�(��A�>�����P?d�B�A/����1;tp���_{d�mݓ� �9xO-��g�cr�x�����ߛ�*	m����x ����'PJ��rʬw���I��K�i\�0��0E\�+K#�ڽ�@6�*�]r�������p�P}��Ԣ��m2-}�ր��&��$
�"\�����熽ټ3Y>�̂4��އb���y��Y��$/�i�ڧ��':� 0��ܼ��,#^[yWl|�;�}������Z٥�%�����L���88:�!��@k8,uG�� �e�m(z�N���BKsz�O�:�����h�����z~ǰ��Z@9�0�T�����[�� 嚍-���#𗌈Vwai$2��HF�+1�������h=�A��X�o#�l��y�d:�r�s��}����(��R4��D��ˤ��'"�c�1S4W��q�wncI�u,av�$��dA�Y��7%�G���H��v�ɝ��~[������M�����ƯO#N�lx=z*UP1����}��`��lF�W�'%����}MW�X&��1���F�[����1���R�]N���FK[8㐯|Z
�OJG�a	4n��$�w&��=����$@4�9�P}�oe���,�V��p_�nC���k%���˹<��e���L��6-�uRL*n��5��7��i+�7����cBY =�ۤ���G��	^��l�7�:����h�Ox���G�E��v�9��w����T�@�bt�P����IO��M�;��>DhLyhYp�T��o�4�����9�d���;�O����k��=�1����@�-������˄$.�u�tՙ�/�r�4;�Ċnq�7Qi�ȝ� J����U`%ǂ���xN?*�[�&v,���8)��S�v@�V�8#2WM�1 ̖T3z�J1�����R՞�o��%7x!(RZAwy�*> �=DN-���C�q{�^��)]8Zg]��=z7��;`�U{� �\b'/�S,Տ�3�gC�NT5(�f�	����0�^n����ЦEM8����e�ivy�l�)�獉��3�qk4�Zs��Ԫo��;k���LH��Iw3:�,tچ��1�������"Џz;�)�ZJUe�nN%�HRO��g����G{G� ��F�CC)d�T�2����Cs��\�m�nL�$ݯ��yN9�K9D��(*[�<�=�, �Q��D=�؎;^�+�:�0�:��_�o6S�@��B>�}���3C� tY�y����^p7���7�t���yؐ�I)��'!�������(���c\;"��:���M	Xy����ܧ���iN���{�iL��Z^���gX���`*D�������lM��o�ު�p��}w�q.�뙏u�*[@�����K�)�1#9zm�O�ZQ2�e�&in��o��R���L���X���(S���g
��鸖#3f��6$@p�(�0Ѭ�i<��2'eR>U�X +��� ���A�ǌ��׉3�`}v�Nģ]
�� i���JN�����e(C�K�o�:�S�Ѱ*:K���G����8��$7�h��#F*`F\{a��������.��U�x(���D�$�9s�n?i�Gx����� ����K�p��_��Ģ���͜��?j�б��5�i���+��Gܒ6����IGQ��$����|��������:�E0B�љ`���BN��R�G�K2���Ah���95}`��am���d�k[��6�Nc$�v���v	Q,��v��$S#ɭ�}��z��W�����D � 7/�����^�<�P�7��t�X8���M�b�3wC��{�8Q�I���z(wG��m+��Vk�^�-)VS�}d��\��4~���#�-F�G�F��%����EN�\}DA��X�~�=8T_�	%ܯ���|��4s>���r��%��h��\ҽ&�y4��V����Ą;1h��Cvf���1Z��kw�	2�m����!��������n8�C���l����VM����!��<�Vkİ0�D0�!��Z��J������NQ��a����p���կ��?'J!>��%�l�):���M�����2`�屲~�@�r(�xcj��l��=����{c(�L�^(}Z���ͬ�
PW���^��������K)��t�qv�9P�V,��@��Lw���X[?���j�z@R����|6ay��{K���-G�Y�9�3��FS+��<�?vH���V�*4Bg�q�է����ؚ$#�5���f�d�a'�$d�)�W@��<�-��cTr������̃�i�� ����#�w3h \������!n}T.���߾���\.���rU��I��|��h�����Ř�rǵ�d7�����9�tO���b��*4� ߿�Ⱓ�3$[\���ّ\�&ղO?v2}R�$;�?��Q��H"��q5z�/t��ԂY(y���Tc��R`}��Ǹ�d]��Y j�I�x�L��l0_ۜ�uE������(ˈ*�'jK��q�C��^��'�!�s��q�gY)���V<d�RM��K�$b�6"Ċ�#_�Z�OF?D��yNc⢭���e�Z�ty�G��? ��'jx�iޒ¹@�ҹ�˶�R2��sm�k��uk,�)�G��'��x����:l>��
��4 �c���Z?礷�!��W?���C��r������־�%/ı��u|��	\J� �0,���Hcc=���a��Q?}i�@@�x&��/+�̑��kq6K�wB�S�j�$�s�&&�/��sl���v�����W��7�	>�AP�,S\D�;�R���n/ ;f?�!��+��GS��bȰ�4�������d%q�cΝ���������ow�;������I�5��p&j
/�RĂV�)���0wŁ��4�XxR�CH���$(�h,pFe���՚�0�:�W��Sg�}��7*�uTY�WXg+�Q[��-h|L��~����l׬�#�m6R^�^�/4s0��8��*-&eu�}��Җ�I�6���7�F$��.�	<W�1�w�Lv�ȏ%g���=�why��ߒ+ʫ�xUh��i�J��a[��`�{��)�o#^t�uv������ 9�I����	�VX*��0Պ���l[�`=�s�;(�1
�m'^5�	BƘ��o|�ra��(3W��~\��,���tӲ^dI	�M�pK^�R{��s�W�\3"=[�����<:����(�[#P�r5��'A��\�۞��QX�ߣҼ����V������ET�$1(��	����ΚR�K��3�a��>?���>����}6�з�
J͇h�����ӺQ�TJ���]��*\-V"���[W�Z23ҳGֵ��[�Y	#Q)��|K<�]aU���`�p����f�\A�,بR��̏��\L:����R����^���I(�A6r4/�[����6�!�>�S(������$^#Q��S7�\Cy8H�#���C�zU)I���p�=4��.$����6���X%~��:����xf�9N��¸X�(8�F�q1�M
)�W����}G�
[�R��S*hŀ����惒���s���Te$W�q���>Uw"�O/��~�O�����5>Z:������e���7B �TP�sO�X�<k��g�j �)��W�p�),:�l^��a"$�Rdzh urΗ6WW PS5��m��[�&��t$k��)�nCr���`�������U,��N��R8}�Ʃ�N�s[5�����*_B̠
ȴ���x���ao���M|�%�\�Xc@��D��Y�Y,ذ�|`E}7z���A���|���Я�G�xSL������,�e��u�>��E�+0�]�RU�{�-ǻ�v�N{���]*�_f(,K��%Ѯ�^���K@�b���y��ӭ�)�ۯF�G�z<�]�����>W��m�!6���A&�lJ�y!�s�"�m[G	7��ޓ���n���h�b�����	���Y�ǟ����|��2$Ef)%j`��l|2�����!�
EV��!h�D3��2�;��ɪŜQHJU��Ւ�o�|Q�i>����d����h�5d�{�<�Ex)�K`��g��g�x�Q�7��_5��8;ey��z-,5M�r]y {u�S}u���&��&�@��GlAaY���� ��c&��5M"�"x4w����7�����\��'��EBҬ�����bOBw�KC��x��I��D����X�q�U1�nݦt��p5���e�]�Ԍ �So9+��whT:�Q�������=�S��k7�*�"L�FH[�g3�E�l&��L_���co�~4�D����B�i�Q����F��(�ybug��E��S��%�����y�医s����[Jk��Sj�_G��=+|�Ƅ�m+���Y��bdՏKk�^K֬�=TsI��zl$����r����_u$ym����4�=xQN�v!2��*��\K��Ƭ<�U�!�IKO�rX�{0�i`��Y1�O:Ff����mi��j��_��&�	ϳJ�6�o(�!0���$ ��=!�铠GӜeό�g�ѻ_A�v�lE��e���0�%L�I��A���Y������rl(TN�R�����݆�u-�(`�����0���DD��K��1��6�A���F��5�c#�7��U��)��|�N��hTc��"�'�C}���K�R���m���S�v���}�� /"y]n9.G/�p��R���sz��S���k.���5���-�Vv�}oU��=բ5m��[��3�0Li���:%�][�\*<X�B�E����U�)��y���\Y�R.��������ζ��ܻ�^�4�%���2�h���HW]C/�k�{Y�[{�!�K|wGt`p�,g#�V��GΆ��+>���p�H�X�E�k��%�AP�����u�n��6�V�0&�џ9>��+5BR���"�`}O}�C�n�ShJx�a�4�j����+�v�|��N�	7�܂�.)8�i��7��ze�r������1\�b��.(���!=��|�g�k�L��U����s�����;�c/W��='����I�i�޺ӰΥ3�(�"sM�(Gc��,�{�@�z.,>��׸�P����v�Ð�_�'M�~�28�#��L1~�]ś2���78)�( �'�܌C��X�pK'g⹈�ɺ�Lg��l[���R��ݰ�n��Vf��ē�+��ƱQF ��r�-�y�nf��u_s�4Fߜ�b�S����5+%��7�A�}�	��>��,*�IjÜ5IrM��ӹ�
]�2~�w�5I���кj�Q_U����hSsG[5�q!�VEх�>8�\��؀aAC򓫚���n��5�:� ��ׯ���gM4�+��9�@b(O�W_C�'��z�p��/)��J� ��f����8����ԥA�R�KK9��a"w�ٝ{χ�,����i�Ӱ�u���:�w��[��a�SJ���L10��5N�Y��j�Y *=K�	�X����G�.,�U�*� ��_��|ǇL�#t|N]9tH
�vn������5�u�ܔ;������yŜ����5ښ�B@qP�[�d��8g�ievbCs\�'P�nX&��+Oe5�Q�ܩ\.��|���+��z���X��N���y�CN��Z�-�$&��fw|�nD�}G�Q�{hs�%�N`]i�Q6��sC ��>������@w�#�)�SmZ82���U=�ثhE�U9
�,�x���I��i��
�8� ?�L�P��S�}��Y�D.��8⸪B%wyj˟1)�m�>4���7�a�k���ٺ[��1�`���c�����C�G`���-��7�����;�`q`��r���Hp\��p4��Z��X.#�"��U2����"�qA�׶o	�ϒ��D�mxZ#�ύ��/���O����K�í���a7
w��M+�SV�BT)�ߞ�L\���Д-�����6��>��FC�i��xfv��TlT��j�V$�v�rxW�$&��f�r8���~j�HR�5�!�Vz|�M��� ��xd|&W�{$\R7�;	�rH��Rσ�졨�ѿoW}��9F1�$;隚}��JzN��\�UY+������s�����LUB�!Ơ�鵞Qْ���^P�7���.B$^��_���q���p!��W8�یo�~��6 
j��� �'RQ���W��:�R-�$����>��v�kj�6x�n���A`<5T��W#)�oq��BG���t_���y&�C���H��N3��ȵ*�{a��񻢸L�1���D��rx�������ےS���'������6H5��5懅t�]ɍ����;��݂@�dE��|	���eG�͋�P�}j!���K�1�nc'��rft��2e�����7�P�iHrɛ�oX��+�7���6�F꘼�w�Аy� 8����P(�-��b3���� T�h)���f��D�e��u�[j=���寐��BJ����\��K�����N;�Q��]�bo�I�^~�2�r52~8�����(�VPi�}k��GR�Ab�/�Lq�5䁥�4Ұ��G0hZ�=j���7lup�����]d4i�m�>m �J��hJ�<�(��̬s�����\�n���n��Yrq�h�x��gz�i��N��Ƅ=/>�늬�]��jE��p/?����4�Q��Jk���W��4���g�5rxl�S��=�TA��6�x�H2�d󮇓�IC.R�\���q���<=���^f�=��4aN�˵S4���-O��/R@}/� ��'�j`">��z�&ਬy|{D��-�$���ɠ� =�N�Q��Z��$~�7�g)��kP��M�y����\q0Y��M?�#�$���u��!<�g�)
��.��	O�Wj�E�*�&*x��Kk����j�|վr������I=��:�sC���\-�u �g�#�!̈́h[-�C�����%$|��;�M�T2S� bn't-���Y|���Jl��.h�mF�`�0�i�\�ie,�{Dx�ו�\g4��oVףx-���\b���iź��n�t���ڲE'�|��Pw��}bc�C��6DW-�h��tZ�8k�x��@P3\ C8%(t�D�� ySް���������T6|ت !��g��u��hs��J;���Ї�.��sI�TD��@��E��`�	�%��L��Ӫ���ں��i)��i���E �A4<2�>��g����C�d����=80�|���U���#0.0���0֔�#7�LM�f��t���`(P��_uw��Y �vp�R]�T�����wFyr�a�����L��( �'L��?C��}���g����D]����#*q��b��;�N%T�H��w�m��>أ�޻��Vb�5݋�五����1ZWmNxG[K\�t��1=n����^i}yQ��v�W��y�o�{ t�����Ⱦ�˴���d�*|��e�^��k�D��%I���k�T`���e������n$L?�Oԁ�[�C��<ȣ���*t!�)�P��{��vi�eY�?�k�Yh˛��$3�<�V��#�8�d�}�X���\�4�q��q��}����?W���3*mn�� n;#��F�=����[o��+�.Ey�8�Ȟ��A�D�7�9b!��5��g����[����ji�hh(t����<v�g�n���Ã�g�:�=�u����T�\�Jm�(�^�b}g�,�a��zs��k��pD�9ot�7�uF��"/���>�*�+Xh��A�)fha�_+�����m[�:�S�hC�T6@��~��F���@rBS׼+=���xw��d`�Ky���q�t�ts�{l�����Jp�x����S=)%�{oKZى� ���N0�(�3���:�5��2�?wB��j�4�<���ץk� �yV>C4����ʟ�=T]5��f`������}�<�T���ʈ��P#���WUA�)�B��c�м����H�k-��xb�!��A��F^>dL��gt)S�����r��F�6g.�W���k���va4��`b�Cv�Q^��;EI���'tRP���oA����?�'�}�t����� �^���4Sޚ���o�QOn��7�z⋝��.L�������E���=��\ļE9�q�卉#zdĖ���h72�x�g*��� qPO踀��JǨA���D�����9�-�b��T�*�x�<~��/�\�&�`�y�%q2�*X�j>2�($�^G�Ņv1�_��L�7b��#��";�g<�9_�"�KCx�Q��T�a�vس�\`�2�e�Z9{��-��q�cZ[���OD\�A��8`KD�||*��&2��`��� ~`I�?d%�+o�/n��[���~��B��_B��\m���U��+T��Y� ˾�.�p����uUf�ZB�Db, r�l��q.��~s��K���@��(��Cݪ��� ���ɑ�(@�ߨg��m������Y��:��� <?�2NI��fc���bԸ#D^�1�G��:8���&>Ryy��Q쌏��;���
;#���B�7��B���v�c�j|Xa���z�6PGN[���a��Dp_��2�����5�0�ٗ�2u�v�lJJ;\�P�}g�[5d1������R<��C��4���X���O8W�T8��&�Q�w/�!Ӭ��E]�~�ڍ�
cEGg���r)����ŀb�?A�¡�������o����lKi�����v�>�3���[8?|)�E�;��i I��i���o�vJ���G��!�7D�(:�����np��":_G2��!���0q��1���ad(���f0�Y��#� أ�J�,�땽�+J�|���P�/�~�h��	�c���`̝�Y\E�h<��EcvLAKBP���P��M��u�\͑��X
���Q�p#�|gSl���{mE**yg�h�0����*P�Q�=�Y���cY�<fl�aO�]~~ˣ2A\�4X3���m皔J�ng�t�k�V}�?��;�ǜ�zI��ўg�}�uUN�+F rh��'Ld���gd�I0�aDv�4�J ���������������ˮ���?>��R��S�(/Q*\x�v�O��n_��PT��gdUM5Ƹ���˲�5��9�p�ik�Z�[�'�
�Л"�R(`LL�����sI�i��-��=jM�L�_BM����Fc[��M5U�
$���*��Ą̺���_�ՐM����C�S�]���(>1.pp��3P��OO4��k�ex��x����T7�^5���4��c!/����qc��h9�Үj%� PP�Q��ؠ�#���*��S�Z�E#q�2E�9�H�4�V��?�B�d�r�U�����R���#٪���p+}3��5@��=��[W�e.�tnI��W���7|~��W��_�4�PB���(U�=ö^6I�";AW�;i`�H1ح.َ̜��Fө�e�.xd���+����c��t\��{j�[3O�9u�b���e�h�.mqU�V6���4Sh���9�G�sb��M:���d��� �W�v�e6~$#Za!1?�]O�)K�GZ���@^o�|����Q��͛�}P9����d�tz����Pc���,\%���*=8UH��шX�T���7������u�v��0�����	��uiGu9�6@'�N/�A�P�Ԃ`7� �x�� ��e�!�gc�A�ĺD���榈ВT'���u�	��T��W#�B��'g:2	 �f�"��RL��-�Q��Z��T�=���3�6J�R�s����T���î�H[�i�<�"TzU����ْ�.��k�	��0��q#��aª%_�Aܪ\b떚jy9:���t2h%�]h��8͠��*�	��{s��'���V�YÊ��#D�}E1�r��t>$*wtr3���T"4�7��c �SBK����z�Y`��>��_��!i�	��s��XZĶ��c��V�A^/�g���vfϤH��^_�:K�w�+:�v�Յ�@�c��,��[�I5�}��r������_��ޒ��A�%u��%iǗ�#���1~r3���}*��}
��:fag�R��ɢ��C$���i���|����#��;�r�y��m7.>�$��+9��P�^!*R�O��A)(j������qx_�����\UgH'�EԦ�kV�A�����	7]���=z��Q���4����*�#T%\����4plj��(+jr��Qh��vҌ�Ś��6�����t/�#�u9(,�g���B1�د�w���y0�	]TD�7���Tj9�X���)���M�]Q�v�A��su,=���Bζ''���x~=�<���ٺ|O4#$'|�a�	�ȷJ�ZZp��;˪~����
q8;�q��]�R��e	�%��s'/\s�y����z��;Up�
-�a�y $�Q�p���qX�b�탥},�<-$r[2k����0�e�_�z_��S��OQ���JnV�cos�"�rz'aV�b+���
�#�޶�f�����60�0Ⱦ���{���T�
J9�܎��S�@N������1!��^T��H�p��[l�|T>��a���X!@B�"�C�MТ?�|4�M��� ���z�H�tp�@'��DP@�]��{Ө�; 1����v?	��v
s����H��#M^,�Ӹ$@��+��6�.	����c��J�k���N��
���� 勃�3��f<��~C�1����v.�F�jK�����t�(�ݬ^�Yk������
��O	@ưv�E�!-]�J:/�M1洃��������\lURd��(]� �WK�uɌu��{`a�g3��9�ԫ�����x<Lۦ��[$<��u�����G��� �%K�j���K�����5 &�u�`��w�.z��`�;{�����d��BӅ���A� }'Z��ñ����LP�/u�� �կ���}�k֑�ӺN��+������]i��s����ՙ�~�	������-���y'��ԣ�hHOV�m�H	���-�rwS��6��9T��K*w* %�l=)G%�M��cӍz%�`��§V����s߅T��,�	xM �˘d�Se�{�̃�N�" ��a-�lOe?��v">g�
 �=^�Y1���J�
����BP���"8�R�e�vX��z�r�/XT�N����iWｮ�F�K �{πz��P����ܢt�^�Rox)7@�^�8�'k9/N�5[�6�3�l/W?.\�,�!5!��&�&0���aYw�)�2�?������xypo[_��Q�2�<{u�<���Jy'��fW��k��5st��̈́���I����9�=d�����G��k�t�јO.����A�̥�����)����K�!h�*�d#��:�Bʯ����3�WD��4�Z"���F���/������ē�o�����DX�����(<i+��2:�8��{AH��|���C�]v�u���W�U(��.G�� ���C���A�!	.k��:�����e�� .w��mʟG����V2�o+�hY�m��^w#�o�D���V_X{��/Kh#{�)�}�����֘cl�7|`S�,�(Qa��˥10�i��\�3���+�k�4(L��J�=��k�0U�=�c
X��BS<�lq�&Tq�2�=ڲ�6pw����x]��#��0}4[��{��k�Zd8R�vwtS�ͩ���i� �����t(�W�n�5��x�if=?D�-��uߏEv��k�ĭ�Qr�r@�/!:^���@��Y$�7-��\��:맇~wZ�l`�&)V��J�s}4�*��V$cJ���uk�O�y�l���s��k�$,ר~�*=� Rsޕ��#C�̹oӮc�a��k%�/��Y��ͪ�K#�O`'R���M|���Z�,t�_����9t�;{�*$��\�E[zf��1-�������)C�����j�:�����-��v��"�UP�P�|����ɾ��d��E�JL�i���B��Rmam<�՝��-S�d(�r�ҩү�|�$��������+�&'N�E%a�ѯN��fX��)���YrF���h��~D���ބL۷X�l����/W�D��&����^�X��a�hĿ�(��?:M�R�+
@�sR�sb[�!��������F�
�&��o!R��?�@�p���ɹ�x�\6��#����9#�M��2�0��1��z�|������X�8۔�<�.��ǆ�0�J���	f��b=q�s��"�䇵6��������$�EF�c3���Yu��y6��$��ԭ�X�k�B �*R%�(k$�L�F7�u�y�p�f�jV"�K�[>�.y��&e�k�#�b��$�ά�Tl;>w]�?PWf�������@���RZ�Y����L;�A�S�ϝ��LF�3$#�N��: �����k\d>r*_�x��A�Da�Q�W�����������Ф�\��9�C��@
%��#��F�U���CA�Ƭ���?Z�v%�?zy�*�����"Z;-�kh�����|��ΙxT)�����Qâ��'��k�]��p��� ֆ[,�C��9�~L�a{�{3����XQK�-紼H�����c��W����U2�	a��ht%��b@n�~{���ْ͂z��E���	#�q���>������^�Jp���Z#�g��դN��i�	Ɠth� 4��@5+P�im/'0��I\y��.+o� t&�'�N��BlN��B#w*j�QU����$]��nȣrN�ו�1mHOU����B����Kd4��
���@52k��6���^֛�Y�L--�[o�SF�
�F@�h+8đ�!��0��Є���&+%D�8�׷@�.����t]�o5�J�����;ס�+��D,��eG�h~&8 ��"����;�J�Z�~�[�1�h����)0[w��{q1��:�,4�S\1�L�#���g�v<O�\�M�qr~�#��:���t*���ʬ1���7藍�{���X���HbZtpc�K���Bo}�]OD[�&����"m�Z�"��ю��5E ��[���G.,��̘�k�;Nv�����°���+�D��p۰��Ν�mКyg����Hg�u<���7��%�W��إnt���Y�M���g��O�ͬ1�B�5Ө/�bl����TMd�(����&tk|�v4�����]����I�� ^�;�͈]����fn�d��1�M�x��z�T5_�*�4��N�0[���6�໣B|hⷲ\��QY�;;֦L�5����Q����9!� ̕	�<J�d�;�=�����ÄH�(�8]h{V�1�e�%�A@8�=r/�=�<��� H�]]4n��d?�T�>g:sQ$��tf�T�%�F+ǻ�����ka쥱,�����z?*�X�#���܀��B��/�@� �����G��DWa��߿��T�0~[��P�~�9b��`j��j��7Z0�XU���XG;�i'�g5��+g���rYj�S\2^�? љ&i�ƽ��ai�����g�'-���_�$�A�'E�E�
W)P�$U�`"m桦o���V��9���	FRD+�:`�;�~�3P���Q��׈��V��Z!h%��f��/A�PbA������_���ǜ�mx]?|j�p:
��@���}h�˟�C� ��L��?�ۈ���;�/�R)q�qkP(��Sw̞�'$>��d�{-�8���g���0o���� (}3G]y%�����EHZ"-��3>�K �G���]�lU�{�ɑ��k�>����8�NjPb�NwVK�ݑ�)B�$=ȕ��􉜐,}�%u�&힏�"7�p��b�d&�\l��"!Q���c���d 1�՚�|�"���F�Fd������8�+NTPEv����
!�ԥ�Eb��xe��;	�qc��n�O��+hȉ܌5�����;{d
�s��b����O92��i�8�ĭjڻ�P�by��qVIik�����#���΢P������ڵ.�w6�L���s�hm4����.^o�D��J�֝i�z�U������?��폔�5޵f��E�PT
k#J��M�#�R֦0H(FՈ�W=3�/�$ɲKe�@*�3� �h�$�X��D�'7R�DK�xJ�?f�j�?��q��wh[rbb�a�Q��wu���#�2�C����<�9�;�sY�'m��'�a��G?�l�3i��f��IF��I�q�3 ��/P�;�@�k 3װ�V��=S�.
f�2��S@���X&�F�s�5��B`,���L�1#�jb�m�����X�]�����M�X�Qv��Rt��e�����N��lw�v.^�����56�l[����� E��Z�aMMOE8Y��������td(k�D�����F�Ф�5׵J� ����(�4g��_���GGZ}:{o��H��� ��zWOq^6���ơ�O����﯁~�_x�I#���E[� r,.������D/z����Xx�w�G�,�����Ic�S�Պ���TZXث�#�f�C�t�ܜ��r�j/�^����y�F�Bgl�G�H��=��_�h���$�7��RQ��b�p����hgZ�T���]�YAk����l�3�r��C�>�н�l�7Ś32F#�6�zS1�0n�_Ы�)�N��A�x�=˕F�u��ja]#������D�m��~E���>NN�� �+�,�_�q�T���?J�^�� h���H�sT<ơA���=B��yh��l�v�[�����ݠ�����6vm�ꕼɯ�*ɱɈѴ �D�QQ�!QyC��&yng����7L���cɚ0ZϞ���BZ��u�衙��h,�^�/W���� �E-��L�����x�G��x�ƣ��0O$���.vx��8=���J˜C��8�7�A�Z��x6|�������K�R-.�H��dM\�s�h��@R4H���3�~�t+�vKE��M{�X�A���b@2��x���٬�\�V��= �b�ɱɼ�����]_t�l
��L��^uEºGVC2��ȷ��O`�7�8NG<;�o;8�����IS��h�\��ãAV����[�!	Obb�n�k˪f�ȉ�Kx?��z��P��?�_���L��]4'q� ��/!�&.����)k �EdXq�K;���n��p���0��p6*W����p����w:���2�"l���y�JbM\k@U0�5d��@X��c]����e����#���O^y���wc�}~(��q��V�@=Z���T�,����.�dL�SDĆ̌g�أ78��+�� ����E�s��+J��r̓to�� I�E�V�n��|�)A�敇���)[f8��eFP�#�u�պ���R�[ޤ5��敩�c"��'�2�p����щ֔Y��F��5ՉZ���;ɉ�{ƷYO,��f)/Ŭ3���p���UMm�(���
cU��'A+�����-��3��w��Q4O��g�	�L̉'ѭ��!W8���0W7�IZ�78Mz5�?뢆4�H���㻄�{o���L��=ׁ����&^q�|R��h�F#sk��k>c��B@�R�w�[Q��!�O<<z'G�@/i��Q�I�e:�N��+/��?G�Fhqu9Tl���$$ �
����Zz��������&3��qߗ�ti���$8)w�׸��J�C��O�P��a����eouf�f��%C�E&�m3��~'$S�Jy� �_�q��zة��u�~2�9��s;S��T;'z����ڟ�˷��j�`9��ƸX/�����:Vh������|��1�T��yj`�n��e&(Ǖ�vs���wɟ�3H�m��y�*	T�佽�3-~��>Ih�/�� �}��xzA�ɺ>���6�X�o���ҿ2	2w.��5u(�<����@B3���r�>��p�Qy�г���b�D��>��.C$=��U$'��+�$��9�'K��J ���%	�3pg~Ș�$��4�׶Z�G����x��螻A�N�N�o��xz<�gi��<������I��nƥ��s~L���W� ��X}?tr�����Z�}?�W�8D7�x��
t�m%��[iy���x�>���ㆵ�;�Ć��7FA���w��/ĕ�س��Z@G�C肻/Qb��$"��ˁ�j�%;
G�\��U�;4W�����X��v�.��yyd����PM&SY9k���@�?�}bf�h���Шu�7w6��u	�NªuR���'$yU���-Ą���R����0w��g_��3�����=1$�R�m�߯��$�:�-x�m�ӛ(�V�f2��q��=v���@¥d�/R�:���T�JN2e�}���C���(�~��������F�5�xCEi �e�=�Y:��L5Rǉ�@����9|������ه���L-�-+âP3�f��>���;���>�
LY��<[�˲(ՊeMTR��,�~�"��\$>^����Snm8ߑL����Y���k���_��h���d~h�R2�O�C��otK��	72��'�d.;�3e�O%vD��M����kI��2�bY'r.O
w8ärf�f/�](/'��P���Md����a��LS��EZzLJ4^Q����� |��]F�*S�\b�@��*��>O�CG��{Z��J�h ����N_,4&F(��T$-��:f{��H޻�x��?>DV���vaoY�r^J?I�3���Zl�L:�^)ö R=!\�n�p�H����:S��[����8Y�
O�.'�7QPϹ����qz��4��U_}��s�1�[h����v��K��T����%��|�qM<�k��]w�M �!f��B��� ��u,����_hD�����-�t�^�NNE�%7�Y!����p<�nMdV��$�8��?c/Io�ҳ��������T�ٵmM�^B�bho���iSx^��f�N�K-a�\D��#x�J.&��Sܭ�v�C�ݧD�@��ǂ��6pT�4��aH-�h�%� ��xH[�5gh@��6Yu���"��� [pl��y����ď�^�T��fw��Q�ƒj~�'��8D�x����d��`��ƨb��k*�s��)�_�ZBM'�`$|x_���x����z=Xfh��Ѯ��1~R�ց�&~=��8�$觗���|8��G�<t}�����,���-K���5�\Y�8B�C�x�O��PJ���
��[�xX�N`��O#'?�o�Ӂy5�����&G��.7�\��S�%���%xup����,�o\���Bݡ��إk�����I�R�z�[�w�*X�f�]��6�|���H`+���0o����h�B���̞������'Q�W�5�P9��v7nkpdR��	��ykwF �y�ʁ�[�_��u�5<g���! [)�:�Qp-,a��Zb5��7�; 6����;�^���!4�o���p-,��Ʒ�}�g���P�E����-�����xx��#�Z�EY7�:Z�M���1h@� D�N����J�Ȥ�u�˛�Q�8͐�6Ki��5� "�� �(�1�%����H�����dU����(��-C-�凲A)�_���1O�׭���p��Iv�W.R���3���l��T�5��:�5^=�Y���S?��
s&�l"�F��Ic|$g�H�˭n��
�����@g~��;�M " ���ރ83{�PJ� ��+�z?�>��+��Y�N3�#����H�i�*O�S&���<.O�2��U./ޮeʢ��Tc�QK���,���%V� ���X����DcZ���%F�7���뀆��p��%ԋ�VW����l?�!��z�e`G��E/�<���9[F%i�ү�ɤ�sv����@��G6z
��}���3���.,���J�E�q��v�=�6�ѭ3�g����>��%�zJ=��K�)(6Dr��-���y.M,�I�����7�v$^d��Ӗ
��b�>�y�AA��*W"��f��Цf��bM��#�Y�x
Uy	Ze�hgd���݆�Z~�ゴ�V��/p�~o�5��ɹS\'�����I��z����	�:��p�o��{z]$����1�T3���f�D��,�W](�9q�5ų�^��Xo�#��|�ܔ�'�1�s�I4q�բ������?	��o`V��� #��$�[6��a'��<���c��7a��U��Լ�A�H������uZ+�nF9!B�����n��R7;ۻ�4[N9��6���@{�d2j3Jw8��l2�a���c|��|��z�rw|�-J������-�x�Ps�����'�խ�� �L�#��|]Ha��m��T[d�7��*es�$Kݝ"U2n����)�61w�8�h�'��Q���UFf)H��m����X�rP7� ���<���&� ��O�����<1odQ���}�VOR7��f'����{���?�3s�t�Uk�����6H<7�~�@ýG������dt*bN��ub��D!�~P;f�r����!?�f�A�����띠��8 Uk� ��*�H���5!��S�ԨW�S��c
5�*��j7�ü�F��q��'0e�.^�����ӣ9�)�=Ąs�G���N��6� 2v��xo����C�Q���֦HR����z�Hc���:;�;х6T��I�� 8��W�uS�W!6M�N���.��HX��A���B��6�zs���������nw���*{qC'{:ȑ,�/�k�+B!��^����P&�N_���RY��M�lΦ�X�*�d@k%J�N���w�J漱Pzi}�//���۽.$e��O�ia~�Ƚ����R���h�<��BL��?5�91"gto	t����C��0R�de�B�`'r�'�����x�Hk>xn1���a�0c=BI��1���#��T�y�Y��i
-�nl�(Z��s)��ޡ�1I�"��~ZB�Ӌ�3
�[|�?��.��M_�"H#c*�4��G��=��.B�w[�s�QEسn/ȓ�Oi�e`	3��H�c"�4GoiËzl�Ds�K��.���0�Kԁ���L>޿%�y�8�k5����������:���2���ڛ��T��b9a�^w��j�f�J}�R��7�}��ߑ��c��L%U�����xA{f��X)������NU3D���/�	���k�����p��c�~#��N�@�����xA��0�~N���NQ̾\\�#َ��+y3r�Wdv��C�oZ���^Q��y���:���B�<	0L|/��Y�,j����dx�oLj����PI�(�n��`�z%�d�@��E��r�-pӚ��d���������6u�Rn�� /��RA�n=�Y��B�������S�7�pn���P:���-���=�Y�p�t�ƔT���;��v;9�眭��3l�F-`F8���f<��lW��Zi�^Iݴ�4G�c�6x�eB/�1Fh��wS��Q���7?!�Y�
�#O��D�\��ٳ;x��>,�I�ZV����=���x�����ɽj�t���vO�������������ⴝKu0S_�א��+���� �{mjBY�IeU�+%Rp���^R�$�v��o�?���wP'��������Pdo�/�h���J�)b��}�5��_^�vG�;�WhX�2Oa��\�H�D��5ib���X�Ic4,�k�=�xe��&z�^�*sq�h}߅���Ν��qx���d\��֋��'R���P�$�`x�|=/��6�3 �]I��H��5�F�3�������3ڌ^M�a�� ��A)�"���dS.�JG#D�wz��@��#.|�qHB*��0�� �t%�P��x���zG<B�]Sk�;���cNe��9�t�fح���;�y����k�7d�{M0S�f���T	Ƽ�L@�IGo٦R�K{(Z�~�B����?-�K�Vn��G�8�!�h�O����q^�ޖ�����C��޻��~�+dJ���6Iq,m��K�y�Y�S0,ۤm���Zg�R;�,�M�wcG���S��H���碲�*�=)]�60Z*��>&*��τչ�t��1!��cKY+ϩ޿~�������~�R�F�-w&�s�j�ћ�>ԟ���N�I�E1BjTI�ѕ}��v�Z����������V!��7O
%������Gcҋ%����������A�X��_�BPZD�HWsN�c��<�!h49�I���,}aL�/˨m�n'��Ƽ�`o|f�N�5���C�yD�]g�g.M�QA�����^'�t��C��^E�[t%�mc����P� �C�IO��'S��w�p�����m�Ox����U�w��%���L�h2&l�}8�ư�ٗ^�4ZP���NN��@��td�i��>\�H�N�f����3�A��'���E���o	��b|�8I7ٿ�ݙ��a�@Ph�t��LFd�y�-�v0�i��8���0u��U��Gd�� G�MF���K�|\���>���ɡ�Gc\t ����N�=�Y�	�34�&3%a�߇_
��N�ʟYe�!a(�fK������<����ǃ)ZN�珧e�X���T� J��Sm(e�Rn��Ϩ�Y�U��B ���µ��]�[F�m5\1B)����,��Ka�%?tڕ+�ȗ_� |�.��l>�v�PD�MN�˘�V��
������z$��[�
wr��f0���b�J��yU:�[&ڵ���ӓ��C��TL�'Wh"-7���)n�!�4ovTQ��.�>Z�^�1����޳�,��lL�ln�G趹1W�(��Cϡ3�7;�^U�ӆ�!�:M�=U��A-m}��Z�Vi; �� �Hn���s�D�̼/L�}�t�>�CM�r�v���%��gQ, ����HNw���cs��bW�)�e�F��l��Ƒ��0�3�
o6�L`1�u�ww�q9PzWL��=���xVwr�j4�OHO�󞆥��SG�6�v��dW0!�*(fR0�8%�"sW�;��.Fz�����B����/20)\m���R)]��e�9�1_CV4
�"13��:a�,���+�Õ��?=F�
Z�32��',D���(�qL��[O���b4�;�g/�҈2�. �5d�_�@Ԇ��a�$
�Q�読��a��iy`�'�b�O�'�Щ4�)�exE��_`p����.臈~��7�lӉ�@V_#d�j����2��jl1�`��W_F��L�6���jM�#F>��ݚ8.��R��-�q��U�����"�\��K�'|&Jނ\q�5f�E�qog�pԡ����K|��Z��?�}�t)ض�2%[K��q����10�IX=_I6���sv؍����r�YU����� k����f�S����K�_�r�Or/G�2��� �A�'d�>�t�q|r�ͧ����)Nn����:���/ԑjc. |��H��_��� �
?f��@����oMf�Nt�Ʌ���^{�xC`���hr�<��G�D�z�a�͒ �6/�0���ku-���g�i�� 2n%�}�a��Z�c�H)�jK�E��3�;"����YW�Ul�i�R�KA�r9��]�=�i�����Jj�oh�a���-�g���+�zh_{��2�ʢ��e#��/qԦ?��ch���՗�x4�n���\z�#�� ��<�KI=��y���B�ٔ*{��D�d��x-���L�
�X3�p?��eɉt�	!%Ͷu��2��FHF�k-e˔�^q+c�Z���:�(�i?��[A���ծ������&�]�63����[<i7kϧ-��]ѰK��:[8=�|���p!�0m$�{'�	А(��A�H*7��C���Eb�D,��L �V��
��@�W�i����!�4 ��䶪e^ ;{��A;ăY�v+�������"���V�s�Ɂ��������'O�-Tv������W�r}�'�ǟot�#����'��������QY�c�ޫ���﫝�#z �G�ׂ<^4E���Cz2DP��ש�}.���=�@o֧��I���5�?V��6z�|��:Ș����3�[�bxg������+i�.Y�
�)w�)h;��
+�8@Y���EnV�u��T`���i�y�s���7Ƣ��3^�hoh���:�`z�=<���e#�(ߴÁ���O��w��ƚ�н�(�禴�C����c�[�W�a���ĻA#�_��j�� S�$��sґ`����U�F�(���ݵ��V�du{�mka01`�1<�O(v䕱l��V�a��ui����<�U�,{(�l��%�z��"����6=-,���/-�q�{��N�A�Ox�h��G�ez�ha߻��Ҫ<��>	xn��=_���I�����DYl��<G� (�~*1��.r*�t�Q���6��c�!�C���2 �k�B`��Q�-�J��Vc��{*��6�}��y`t<N��+��Y(YlM��#�O��{�/�-b�V�a�AG]fc�u�=�w�Q���
v���P-]�a�Bo�|����;%�FgY�)�l��7S@��&M�\�İ�90N�/.¥���r+���e��)��g�d0W��j�}f4�FVb�&�3�����bG.���n�ڨM�g��MyJ-TԖ���0��Ӈ����Ev����y��w��f�ʼ3;<r�eH��{~���
}w+W��N�}��T�v��mGA��Xm8����][�u@��8�ެ�7��w�(��jx��1=,ʽL���2M�����À�Ә�U'rJd��Z�,��o�D�ze�Xv�C�H\Ϙ(ܑbOG�>�B��d�R0ί�@�%�=r9  �[��<d��1�T&[ \����r������	�.����d&\�ؤ#~3M���(���4|����K�y��Lh��?�.�S>y���/*<�^���քu&<R�@��aN�*O�\d[�3��!����{���g�rQ�f�ٹ���?6�B���x�H�V�oƍh��qBR���A���l�#�i!�Zf�ʙD�֗���� �ђ��x������A'���4�̼UVB�,�G�ۆ��	`_�/�Y?OhGJ��'��e�M|�v���4�@�Z�C8�6�.�c�Paa4O"���ߗ�>� �w�Nӧ8,��>څ��#��2��[��%J!�i�q������P�*�)���ԡ��Pk��<�j�� �S��;I�B�еKFg��%d�ƠߺJ�G�uߍLj�!�][���t,��Í_�zZ��	�n�3�P�CM�i�`G��6^�_����xq5ժ5$��u�Vr�T�њ�:-&�OD����܁�/]b�'x�w��X�ND�d�&	��A@m/�#5U"�u'�@ޘ�x� ʋ��WT��-�ﾊԬ����i��ZTQm���[�1�K6�����|W����B|�炭��:����M�e�V��Z8���`�hL6䯈z�H-vd�YӴ�+��X��stT|��l!�623A9-Ԁ�~�� M�rS�{6�iy�����֠b̝�!Ҹ��З���zр�{w�|-W�1I���q�b���|T��u�o3��h[&w�����2��������<CK&�_�җn�^4�c�u�-a�U�:���;⦢�UZ�;/Rt\�$;�9�#Ɖn��l\[~��_�N;{�饯2�Î3�,"�hP�%�"[��MA2M9���Q@��<7i57#2�Z��^�?f����	:���*���>P�S�N�Ecwɭw���fF�L��e��/��4����"�C2�*Z�*�]f�0C ���kt���^f����v��A>�us7(Sv���S�yp�W��W�s����>�i&�`�M�q��ھϐ��U�a�%��<��%N��<��,8�Q�@���c�:ʓ{�">DC�.�@��r�z-ۇ��b4N���zG���>L�vm�*4�LRV��ʛ��O���J�_\T�9��,fu	[�D�j�=@�ʋL�Z!*c)iIN���>��n2��_LʷbsS��uC5��6�Q�����%�(a��Z[f*;[׼���g�f>�k�A^�_$.�Ǣl����a��?l� �9m���N`U*^s���_&뮏�u�>yaڃ٥di���&����@qn9�͗�����h�ax+ͮ?e����ss?3����d�T8�eӶ���+���������>h����Fݨ��{������ð����۔�/��bKB�t���`!S3���n�~������uMo��א���S@����s���2) �s�&s��i��a���0��A8c�ݦ�v�/$
��n�2m�P���D��u�%����U��AiK�2�{ܭ��i�	��jq� ,e�!+�6���x;�>��?)�g+B���.&g�vۊ�bYz(�J��u������dW;��IX�oҿ�0C��N��:}�/TQTӃJr�]����v�?7�ŒM�B �_�0�Xء�Ks�Z}x�s�ˇ�W8ɻ-��{:����ˉd�h����l�na�hԯ�������w��C����p�R��n� ��S/ ^���Ҕ  ��ټW'��	~_�n�l�:�_�[��S.��P��t�c��-�1��@�b@64�j>>�I�z��ևT1sq�6�Z��%��_.��O����ަKR2�-���ٗ)���˙��z"re��eZ�!�:	�Om�MN ���f�.�1����.י���j���2J��j>TL��'�u��W���o��Ԥ�1���E���������(c��oB��l`WVp�=�;����!@�_ՎW�X^|j�{�wC)�������<<���P��'v0�}$�nj����0����&���X9���N�w7�:-��c�����fD���a4Y�3�^��*Qԡ0�jm�u`��� '��:��/a:m\е�K����������U� yF���`����w����~ 2xrZ��!��3��!����˹]�XE-,�-�,�i�j�jkϑ��1���p��X�Ŭ�G�)���V1���DǑ)MKM�����k_��ͯ�`b���ѩ�'M5�X=i6+��K��{��+�.���/�j]��Z�w
`�!�|ӊ�#�m��"{)���vu�X��!9#B�o���O�Psnb
*ww@Q�S���6�*�x��ip��@r�9�EB˂��ˬ��+�d�%�ZN�VVHc�i�[�2QlӴ����:*����8�!��A�Xx=
CoY?��Ժ�]��)4֤��&��,���O�I����Lݾ�a:A�e��K��%��9FδP"�M@��E,*�$l���G@�J�����b	�@�^M���}���~�-���QM#6h�i��G���Zh_��鰋[�ܞ�GИ�W������k��H>��|�A��(����o���*�Gх(�~���i<�a��*�s�D�9���;N�)�h��T@�(R�~�%|�K��l�Q�:�6���;U�5M�������6����מO7��`=��g�(�� ����J��[�Q�^��em�����s�Q�,�z��N�}8.�{ �5��|
 ׆����sۯJ?����{7�@�yx�S�xgM}D!mښ�ط��H-&i�Ś�YĒ��:7��\dF�N�2�vr0�ޒ�`�N�=w�q=�'6y�]W'I��7����n��x��( �vg�8�C䗉���f`:���b�P0N��Q��;iP�w��P���Zb>w��!�Ŷ"Xp/ܛ4�)�RT7�Gr����ڀ�'bʙ��)ߥ���>��@:��wc��w�:P��?�Mf������+L�Y��sZsDd��^J���ݓ��6�./��Hd"y�*dNT/*�ϵ�3�ۢ�F?��_8��V�Uyߋ
��Xt��ǐ� (T|
�J/��3tx�e}7K��'��x�f����$5䰫+tA�A�5�>���e0�x����ƑJ�:tK���+�5J��9��x4��,�`���A�D�p_��ϰȍ�?�� M��a�	S��I�84Uz�8��G.2�����IN�;p��Io��\�-�{-e��j�L/(3�7� [r���� ���'��Bf��}o��c���й����A�:�%�%���9�:9��A��s�s�������=I7�IZ\�JU����Z#�uҧ��#���r5nt/�S��a�����[�ԕI�V��^b�'�:4���f��t�_�m��~���^*��W��497�oNjP�(���^EUo��Oj	�/��
��ip5�a%0�g�9j�I|x����"�����	~��\�q]W+m0�7����,0��oc�#�60�-��R�.��ԬϾl#:_�Sus-�?��;�o�(��6��*
�B�}�|����|���0��+t%�Ѫ��"R����k`�̓�Xn��anm�6�m�l9dP���pP�\-�"��J"k����c6Z�����+/eS�~V�����D,>AJp�2<�ٔP��m��� QȠD�����B1odo��۱L���B����Q����;<���Y樷2�����H�*���f^v��	�q�8.�.ǝ!�,��~lcs�{a��8H��d4+)��~��.3���x���������M��e���7F�O�B������>&s���zXWm��qf��b��$�R���.N���s�Q���>������r��O�<�F��k���m�O�*�ʠ
��$`�sn3j�<�5�+��+'�c�~����mW����ǩ��]:���w�cc�00'�EP�|�ьT7`l6��3T�&����Yv��}��j�^k,�;�F�K��ԃ���6J'�~°8��D��P��?"���[��B���q�}牝j�>�R�ܑm"R:˟ �{J:��uDI�ZZ�O '22]<�e���]�G�fC@V�
���	zf�3��j�r�A�	`�Q� ���,䞜�A��|1�Q�k�����^���j��9�r&ըH�q��������X������|��;��B;��Tڮ������P�Vs�Y��cT�:�������E���n[Vw4]�/&���_���;��#���+�
�:�gG�J~@�̒i��Y�`rm�L�@����߯Ь �\¬<@�{B
�t�4�D��H`�\�d���H_x�>�I�eɝ��X6����bLG�	�5�k5[:Y�8� Z$�����Qg떘ʏ��1_�fg*��ַ��+$Z�� ���`T��Ss"Mo�W�M[��1t[����<8n}�+>�x���tr����7��	��-��`'����C�:�y�����ѹ�4
0�^�`E�b�
�k�^%�Y���"�ITiY4��go>�����9~	=\�i8GfΪ�#�S�!�w����'��؇ܞa�h3X��J~� ��%VE�Xo��L����A�i!4�s����љ� ��.@���K��o�N�S�3�1��t�	_b!���@E�K�9W�U���@�W��V.�T:�����4;&��� ��M٢�����5�YWU`�
�z n:��0�+�rȉp)���3��v\���4 ��G��ç*-������t��Y5Z�*��A�)�J�S̿���(W���={̶]�6��32�猑Y�}�������x �~�}!S.Zju+C�Fw����n��EC��u�6E���j*�5��'��3�}Q*���b�1aD/Dd����.�����h�hU(���_r�������������c��؁�==O7
�q��PӁ������}��w'��Z�8�/�{y-�!A���R��ghȢUva���`-���C��Ҷ��(o�����k(��+z�Յ<Aʿ<&�_�ν��Ch>h�PP��hK�9_�]�
c�毵�����ޢ@JK�Z4�6@7���{��,kxݼ�,�(bځ��q�V䫺�#h�������v�^3 %xN���Q�rJ�y��rJ������5��HI����)'Z�X� �Ia�𽫹��Φ���M+�)���!}�e��Ѵ�%�5��* ��p1�ٿu�%()[yf�]Z�HZ�5q��S�3���\K�P8�×ʅg^,���¦�e�5���_�*� ;X�̅K�������2om�߼9>�3`�����;��VG�tZG��;��P�5<���H��,ia��ǃro�OA���Nw�-�m���y����t߭�n�F����=Lp*���.Yv��5�*B�����N�R\��1[X/'	��վ����:y5@�6}|���U��/_z����og�d�$<�kŉ�8��m�J2ZOsWM�� ]�
8ʋ!�0��(�{�\T�R?��`�µ�������Z��`ha�k| ɾG��;x��1#���������+�J��A�É�V��4��D��|:��f����KQS�5��7��ҧ���S>L[�~�9ރsK�CG�ɽ��rt�h+!Π�=�Yj�MНT̫���E^qf�_�ܹ����~$��6��^I�|���l<E�k݀�0�y+�C"��x=Pgퟦ9J�����	h���`�����R§`��m�,��V?��GUVӎ���6X��dsl�tŢ5H��VC���h'OYǠ뉕:D`U�{�6��K�T�	kKY��q��zh�M&�>m$�o�H�b'�|-o5�^3�Vcjj	���t��
�Q�,�v�H���y�^Cۙ��6@�P�X��ܣ�?M�g��8,:��L�[����o�#>� e� ��9 d`�BǏ\��r�UT�?��>�p�0�g;�s�����":������^Ve�Z�ԙ�0Gn�i �#�݅�;I.~&%l�+{y��ymɌ�z#f��X*C��i�l�[�N�jL� =_�q�Ꚃ+:>,$��PJ �����
+���'آ�SO�d�캱v �������&�T�e���y��_m�\pۊۭT��)�e�J�K�.��6���"&8�\��ݍ�֠GD��"Zu00:��҄��wjNX{|��c��,ր �)'L�ͼ��ڤ�*�%���Z�0�vPoO*����)��U���	$[�a�m�6�&�U�?��Ҫ�	�ǘL����D=��#��EPf�ݰY�a�ҫ�#�[[F>]-��]��s����He��I~u�S��m��K�Ϲ�O�0������H?�ɐ�'0��	�ȧ�0�kG
��w�+^����
�1�+�|ʪؠ"�4m�I.V�u��ҁ@d��G��'���������d5�d�8=�N�G̠�����U�I�07��t�S���Ҋ�V�VD*J��-MM� �Ɏ`pi�A�Fu�툓;�Qz<!�q~�$��- Jr���X��ތ�<�Mr�Dg��4�w��b冲,���L,�����r���j��+�}��~��燜�r��\��/�\���$U���):�˵���c�!�H���5BFR�����+u{jr*�a�j}��+GL��Jڦ�N�F9L��8*Q��OJ)��.���Z�����p�-��y��4:�1+�� �T�!�����iO;@�� �$�9Z��Ύ��� FM��~٭��r�愕l����|�������_DQtSu����R
��e�q
w=3 24N��aرs�'�3�0@��+nh��_`zK��,�(�?�����Ȁ�F�߲�Ǝ�bz��C[R�En�b`Q�tP<��̆�bIS� 
M�)z�X��+l˻}�
]�h��~C�i�o�� X�phSh��)����(�V��OKH����Y,27�C7��2�-�vٚ
t�"��I�{�7�_Hƈ�M�B�_՚�3j��Xbg�Z	��?8R�cy�_YP��@	����\?�.Ը��T����&w��veh�A��ln�*5����=˿D��W���:p�a�PQ9�w١�@F��a4Gr�U�lٟ�ZX��.���N
pDm��Q�^��1�o��v����7)�e��Ƥ�,"~
���i�?�%��	jfk�^qtj\�)l`U��B�,{���ҧaJ��ӎep���-�y�y*ɲ���dUp�2ՄX�������m�.w�1��V	6�Κ��x�,,0n��  ���bYĦz��YJ�&�h� ���K�v�\W����<��~�>��m�&tP��FH�ժ��4B�G��d˳+��G���A�h;�mk�&�����V&������}�3�����sv'�%%;��"�r���=\�pm>R��~���3S������5�?$j�z��ezv�6k�垸��*��d���ӕ�qoZ3O�]��#]��N��5 a�چ���$֢@�h1o��k���Z���Vuz)@�D�i��[���v�i���R��c�� ��n̉����M��V��{��+#3��U��g�U���ܺ���L ҿs����e�@�__{m�ڵI4�bTW3z�%盒f��ߴ�d@��u^:�2�R�eF���r���U�圚���B�*��l��"ٳ�l��^�L	\}PK̊�K �@��r�b08,�řilw<Lpg�a��B0�CVL���4�h2&�Y�u�/ �!&0v�~iY�������u;N�A�[�n�B
�$��8���gL��˲͎&`�M��i�b��7S _4�9�ǊQ-�u�u�&H�z2��+�����R-=F6n������F-�U߮��GO��.p#���Ǐ�U�ҐN˷tb�&VG��S��2Z߃�I�F̞�'���I!���\S�<�rj5:�^=��3w� )�3P�3�c��)�^�es"�,b;K�e���~�[��}6Gʰj���bgĸO������#+�.:y���[�������h��~��{�D#�C�'#�שY���x�&ixue�*km���)�$.�NaG�/���[#&�ZM�񍦹h��ᓼO}�!R��,vW��i��
/SF������A;T�bǪ�v�Pg�m�[ya#�-k['w�|�Y�-�X�#a�����H@;�t�E!q�8��2�[Pz������$$�B?K�@�`���y��N{4�97��k�ݙ�Ð͏D�Kh��Fo�H�IL�&���c�q�Ө��29r��)
��Q�
R�'t?�#��!�6�=/���Y�����B��h����N�7�I]�B̐�+�X�H��U���.˨Ůu��_����&���6�a��p�o��J�@��x��z~��N������12��Pd���k�Pic	�/:%��\i��\��7[j`���S>�C�
0�o�V�k�SŞ,�~i�L�#�>[!� N��ֈ?螸3��+>�_�#��1��ނñ����ǚ9�05(�'_�9����+��cg�͌g��KsC��s
�,��M�����pN#ٍ*kT��֛o|��j�D⋄T��P��.4���6\�����#ݺ
�^������'!�{	��ww7�+��q�Q���ՙ��DЌ�v�P@_��$m7uD�_-V��5�ԅ���1�Q���	��t�K�b �K���v���L2m�b&� �3��Ӕ� 7�{~!�?���o�@�o���ڵy�,�|���*��H��'3	�5 v��(�X�Z�����|�b�Κ(G�>�-��u�!�*�y�N����u�<k��T���������F0���6�~E����s�p��B͎{_�)��a!Rֻ�<w��q�d�c8)�h`��9J^a)�pr�L�N���FDj����L�a�xr+�̲{Ů��/π]����g�(C�v��=~ֺw-jS�MG��sJ��[�{F� �,f��^&���V�;�Ӡ�8�f`�z<�P^}����C�����;�&b�j2T�"Q��6[�գp��+ʤ��+}v/"&���{���J[�~��s�C)��޳O<�UĻ5P5V�*t5������_G-�c�N�`�����"p�uA�6�{���IK]�2����ՕW���2�y��p6^�,M�\��o#��H�C��8�$�.��̯-�):'	b���lR$y�k��]l�%�h��H�@�q�&u:�R���DG*�M?ʩ(�@!�� ��������0�T,�yؼh*�Ǉ%�fR&�fo��Z�H�<���@��%������;��4�j���4�����0cb0�2$
�S�l��x��u3&p�E�\g��H���#��'���L�u6Q��fB��(�@<`؅��w2���29�w�nkZ'�Հ�!�!B���V�ƪ��{��ܫ��<{�xƖ�p[�
0��]�u�ٌB��9���Y�S�� ��FK��&�J�
Be[��d*Q��߫F[�@���:o�gL�)�9C=�������d#C��L)Η���mA�wf����o�<M�r.=2��´�	�����`'�!���m꾼�ss����i�dw�% @ݲ��gw���ȹ���5C"$-����F�0�x����AENlJz�ɾ��"�ޔr	��OLC�c����^=-�Ӊ�-���O���K�X��(���hf�!ӻ���_O� ����0�,�^�A�T���9�
r�ikRrA��q��F���ѐ3)h8�x��es�a��w�/g+�;+��W��F-�(6�*�֏�D<D� �<�FL��Os�&�ø�$�������\I+}�f�p^	�j�b��� ����>z�%����f�,�\ �Ԩk��&�k� k�M���d</�&�`�f���'z;oh:R��O���,���JڗVzE\I�<kZ=�4�lǀt�Bw����H�WE@�:�r5��$��l�Z�L|:F�z��ԥ�[�R� DO�,�ހ��\0sܰ.�q�ls�3��*A§|Ľ�h*�a�wne��'a1TfF��g��r(�=F�_]��k�H�n��C@I��u��U�c����$UZ|b����.R��2�k�S�ง	)p��ku}��Szba��{��!:5d�2���6^��l��,�=�g���,����KΑcig�G�LҦ�B='L�W�BS�9�Du��#����4L�^	����%��n�`}co��\�S��&�%�g�֒i�ڻ�V!ֹ)�V	w(�뾡{q~���f����_�t��ҷ��V�X�;�"��2�T�i��;\}mڦ���_����X��Jf�ȏ\�1�Zh#�Y#�o�Lyne��v�[�d�7W��W�]����bp��Ai��ޯ�_�?4�,+��MA�g^
i:湼_@�
�@����d������b-��qG`��n�����&�*��a�1U���̂�y�X��۳��x�6���Wլ�~R$�|�m>��Q�vN9QT ����ItS��O,2R�:Z���ܚ_����m�9{Eݫ3ݹ�F����9v�������"��o�V�8BK���׉���0i&���L�t��4>���j����6���6�:���96�3aw�S.T�_r6Ŀ��5J�9��kŠ��IZ���w}9Z��ށZB����cpNOA�{��Ҙ�tb�֏5!e&መ�|��++�?��јFiC�Y��ο�7\a�78�t�۞Iղ�L�Eҩt�_[��c����|����~\���z�'���&*FU����/��0��tB��{Q-�m^O�����|t���ߣ��C�MTۤ�$���#|���m׫�a"Z�i%��7ׯ���,�|�I_�D�q�uF4}�ز�P޹)׫ه_iYv �W�^Z��=h��B����b�q�]�;����PU��
�9MW��ݱ��s����_B/A(�r��t��dK�Zİ�DL5�/?�P�Ƹ1��]��k���VM�Q=�2ߦ�Qj��(0
�\���|S�i�1���?p�8��T��n���H�kG_���k%�����Y-���U������3�����F�L�^D1�f�f�ClEP�'SAB� �I���rJ	
z5���;q���;Q��H�i�.����_q�1#$�{�H�<{as���!N�'�l�"��ӖE��@R�\2��v\Z��&3L�ͷ����@ �9
Sш5+Z��	>3�������F��#�M��K�y�ض�׭cUJFmȁC=������y/N���<�����m>o�O_ᗳu49�vNO�JN�F��ο�Ip�;S����k�kȔ*S\ P�@B���۟��`֞���<@�,�|'��������c�Ș�����VRm"Ռj�;��ْ5�]H��
F��p���Y<��}����(lc�H�����Īᥕ����������"�XD��i�x�C/b��������UI�	���r?]y�8���#�]۳W#������;���R9��7
*ૂAW�,�m摹 �S:��� �O���۪���]<�	���oJ�1���3SP��D����օ.�,|�8��7e��4,E�pI��e�p1�(���y��\�Z���RJ'�Ox�K�~œ&T��<�7�=1�0�)|'H��l�'�����h�(/��s�|�,۠�;�ӨU	CM C��O��B���%�t�"�˔��B�Č���E�#��G-����-�m����؆���w���[�SF�'@��fĮd���B a?l6�A�_4��n9nT��
ч�nz����|��8���g/����Q���6�����8L4���njh�=�h�^�2ظ_<GZ�Օn���"�p��#�݇��2�w �xw��(Ќq`Tъ弣<!xU��}�J��i���֞a|����@{���\	b���qٝ����!XvRIK�\&��)Y1��cp?n� hv0�.��k���DA�6C���%�оrj&0�m�8F�Ea�C����!~$ ��%��l�"� C��T��ڧl��ۮ��Rs�ʚۢ~_�����T'd�F.��Ն�d�P�4\���<����-w�1yr��$X��<O�GN4���
���@%���q�_�;��5J���u�}�~f		Q���C����ل�����
�?��G��2�Ώ u,S�JT7�E�x��d�ǡ��g��|�w�늞��2��:��#R�_�9+���rFZS���(���+���9�ʎx<��a�YǬb�}z3!��L���q-_�;�,r���ۿ?R�[ao�=pd�3����,W%O���w�w��k����6��EY"������Q91c���I ��Y�F�#�s����� ԙ�6����p����_= �5}g�[k�م�T�7#>�}| +Wm*-�zO$ÓY�+��;s�T��e��
�׌I2�p��BK$�kP�תe?Ǥ'��"ex7�#Q��9��j@�R��O���x)B�%��)�dJ�^V�1��2gtL8��'�
��k�,}5�P����gM��>���JI�ιŵգ��!��4��y�V��d@����wJs�06�HÀ���K����_��Vܭ$n�P�_O��V/�c��:؍�]6h�zh�t�&I�>H!�x[��A���s�A�C�+��6�ז/��c���@AkN�)w��aX)c��Sۆy�p<g}�bR����4��X��t�&�\{q���W�$�����@z�ǽ�f������z�*���n�2����%�(�drq'�fF�/my��X�V@a:S���G�kw�����Mf���-�p_�܄]T۠�7㫢*��h�IiA
�1k���nQˣ�~T�]���N�A�[ٖt�'Gd��*���R���>�RwDv�P�1��xVC��
��,�� ,�u�]�b-V�0���a|pT�97!������+]&j�L��І��L�W�f���\��:�E�3�v_�$�Lߤ�x�Y{$�j��� (#��	@���#ܳ��A�/%A=���H]�i�AZJ�g��V�0$�t��}��J��0��B�������OX�.;��\�e ��e����.Z��-�Ê��A���Bk�0Tփ�ۥS��F���bu:�a'C �,���$A.�L�sj{����;�h���4�:�$6Z�Oi�<�_��k:}]�1?�"L�|.!�c7sG��=oftX��*�Q^(F�r��<�i���<�n�0��̶p��w��#9^�=�c�r0oZ�;��S��Ԩj����s�p`B^��<�'�� �\R'
��׬^�t���%D��L�9vG�;�lIO��´tj(����1D� �%�Y���-�nm�jj��uO���p��F(<6�����CQ>C��7�n�����Ad�][���{4,x��(grE�8|�K{�2��Цi��}�3K��1-@a�����F<ʓ�Еb/��������y��.���?'Vw��1O�.��Q��`>Y��*6����ܦ�K�ĩW9Nt�kz�kS_kt�N�ۄh��!��+/FT����¹��P%����Q{����B�w�Y&X�w~aBC�Xh�D�W>����hw�s��P?��E���4:}��h�طE.Q������c(H0y!q��Wk�gt��7��9���ƍr{f�@-���J� �#�L��y�V�+�E�J��yQ�@��o\�����=�B�O䄀L�^�g#��IpO�]�n�XA���fJ3*J�Ο�r�7�)o�������q{$y��p�IH���
�ʹh���Bb喑�$���TJY=y����r�c3 O'��+��JE�pS����^��/�����C�tvI���z���q�ԡcV�u��$Oͼ�[�!���fllyz���9 nJ
bsHJ3��؊'�ʓ��|%�0?�0���W�:R=��E��T~U�;f$ �U��[g��?��|�~H=�n���Eec��U����c2��"�n�R	IK)$nf#zM�סZ~c8n���c�s:�{}AERg#���c���j�/L���-#�
�-E��4t����7`� �ݪy���Ω#89<j;)Ϸ!.�I��>a���黰-��?S��J1���Ye)}a�Ur���Q�7��-�[�o;
�i�$�䖾!�y���~N�����}��w���?Z���3F��>��(�;mO�v�:�����fp��En�}��/|��������@ٰ̨쉹�����x|x�A����}|aj{3s1�T���/t�zu�i������
��0VCT&F��E��4����(��{���oP^�-M��o�:�g�(��믻��B�JЩ}�R�	�4�Rb���qE4#��
3�	�s��z^�klNS
=����O�R��.{�-L"��ʧ%��-����VK�q��r:z˅y�BBSI
HZe���.
�����������Jح�mJ�Ƹ^�u���4h)$	E��xa��&#�J�iF]�D�˛Qz�RjY����Tޗo��4��,q�`�X36�5q�K�1���e������ �AǱ6��X�Q�)@r�:P�V�`,^=�<��OU��t�����]3�v"x�j����EFU�����F���Q妞{I������(45D�]3"
�X�-�b�RH�:����Mk����ܯ0\�����K��f�x�<$�:`fӧ�'��`eP��8�k��N	5������xP��e�coҙfk-��W]Pa��ZV%*6���X �C�g�i�ď	�j��ٜø���˵�(	h���@���)�0�M�.�k����%���H�^��(7$[�ͻ�_�
�1��,&�9X�P����J��=1�y��p����˃ ��[V�N�2g�����{C ��,6�\��p���H1o ��e���yp�Ǣ<$�Eس7g1��ꪈ쟢,("�p���D!���7:6���IE��I��àk����VF`x�gMD���+}Aoxyc�t[�~�*�5n}��h�9eksI듍iEd�%S,��K^X3�!����F�q0��5=#����}E�x�I�3':ԏ�<���њ�J�� �JįŖ[���ο�̽2I�q6��N���X��^%������ȧmo�5#���u��m@
}g��նc���X�Y?GY� >/��J��t���F,td��J��#�cM�{+9o���c$PC��O��g[���᧏��.��eX��ߍV������V�p���i�CW�`�&[8�H��S$9��d��o�V� 1Pl�Ţ"{�L�$tw囨��zU���α�	����:��k5m�E1é�u��:��C�K#ٝe�R޶S`�2��BI?+�0�m5�wW�C���U�,�3��p<,u��ќ5G8t,�V����'쪕]�m�u����v�U�'��L�Y��::^��S]��,e�*�\�ad�-�ݗw�/��۞�̮��|V�fu��I��k�bu]�=	�-���0C;�ҋ��F:3��nGz=��/��� �R���?S�1�n��[�#������d~����	~�A�:l'�s#s�ŲG#z$:p���g����e{�x7x�wfP"�#�A�a��ݝdv\Z%)R�o8�k�"Xl�l�E��k|���Vȩ�z��?�/t�-1_�k�ģ�]h��_�Xs�?��\���RE�=iO����e�o�\u=J����y(Pظ�>�%�I|�^�r��o��Uꩮ0Q��Uvb�(�;�����*O�1�%E�O�
Qp�>������"�N4*�{+0����)�B��	�������T��}����T��cطi E�k�n�
�~Z���`Q��"e��
:}�lv��H�v����-�%1vU�s��;P4�Z���������3�cwq.�P��#��tӨo(�/�/�K}}�●��Bg-����C�ǔw�� ,���
��mq�=b���Bӛ&�%�[���Y�B+.-��Ƨ{��o�6!�kɜ)�X��q
�2�~N(�e���g�2�È�꯹����>�P
(�i&~-9I��N^���|I�5aG�a��覗)�N$"R8B�Z�Z�Jjq��A�g���u�ƅ�V�� k�٦�wyF�k�b�Q��W��f���8r�8��T�J��i�Y�s>��-/B�Ld#�KL���c�����Ì]�~\-3���W�F�e r(�a���'>��թ �����",��w�����=��S3��j\�Z���2���$�&��,�ҁ����$z������ Nf����K_��ڋ%u���'����)xh$�7�;�~�sxX���ލ��&p�fs��U�ń��cl˚t��a|	�f�뜦
�}2$zEO+f5{��ц˽k�ࣕ�H����+�+��z����.�p��ϋP��au�(�?�rMHP�X@�R6`�]�>�'p���ťq��ح���c�*�������ئ�׉1-N@��NĺT�xմ�o�u�3�Y���M�h��J�5p[Z��3Zs�̊��zj�UL;w�3�I�NaxMc���%�����P�#���;��az�OK��T��{�V�Ul�l�Y�׹M4��^���Z���|����-�qc.�j��$-
�,�����W����P����]!�6,,������ʲ�g����l���.w��S�'�1JΚO�⭊��҅�wJ�\��'� ���\�1�H�m-Ƶw1�r�4"6���I��j�f�촁�8 wv�@� *�p�F(�c�ގ�%"ѿv�(��o�V	g�iLaj�^�D���C��M��%�
٪�w��� �/wH�L̘����g�Cp��j����*j!p�hص���_`�IjM����=�F��9�+=�~��m��:��T[7=����W`!8� 3�̸b�8͜k�+�(-�e��¦���'����&�̇��J�$d��[�U�í��@
���T�6�[W�+\}2��z�q�����b���{�2�R?�*�x��$X:�5&��K��݅PN��f�9�R0�k�{vV=�C��+��5��-z����Ϸ�f�u��Q8��'7۹�;�W���"� o�V�3��$V�HŠ{�2������F:_8�7��pi�?�L��ޅ���h�.��_���Tf�蟈g!�/��/?w�lo�4�8A����5i�&�lx��:��hbLzk����y1m�$!�.��[ԫ@W�{�`���z
3��S|��1�ip�&f�����c⸺��%� ��x��%#l5��~�>�y���bP��0:�8����2A��.?R�h��۽�� "��mmh:c�$�ח���Ֆ�]=\��� 4
�v!F�X��Z�8u+ ��Q�A��Zh��r��@i����,\��|G¼i^��+N�{U����i��a��r�t�����5")���}@M�MG����l;㰙w��������\/�ڂ��^�U�MD�"ǁ�q��$��5*����! ���qVq�ZD���/��ؿ�I�2��#���?F�\Ž�Z�6@�2{�B��ƶm0 �Z)��io�q��9k �s�@n���%�*9��Y��x���	��|�r�m媩bQDSe��tv�+[lfӫ����)T���ڈ)�u_S��G����?��` �
��;�%��yŔ�UV�WXC���{����!C�|���7��F�\����}���%�iQ��c�P<�٪�f���+U`A��0�ȕL@�cq\���5�����&z�:`Q������I�2�r������*��ƻt�x��S�śe�|�e��I� D����4��:2B8����QH� O���C��@�MO�3����֨�Л�}�n�[����@a��޹�3Y@�ݴ�_*~I
���G-S�jP]eg@�L�Ɣ]H������.M�	�K����Ư��F`�б:�&�8�|�K7�h�2��1�c�rC���\oZ,&㹾�YD�Nz����etշKr]֥��B�?t�ݫ�m��<��o�i<�14z�ĝ�Ĥ�Z�������E(�$
Q�Qs�G)Y��K��d��MS����5E+�(*+��8�3vg�V�(4�Ӹkz�a�qV���Qd ��R�ÆnS�	��"�Zq]��*��.��)����f�����١+�D�U?���*b���!�b-�~�5`���_�H��h2�ИY�+N�~4PjJ�i�0�H���G�E��[� ����UJ��>K	'T���������Է��7��8u�x����&��*<]:kS9}��rz@�'FDS�.8&:;9�-�J��?���[�� ۳͛^�?�%��J�(c���p#����6��F�?�גV1����tȷ��]�境�:B	k��u��u��,
�;Ox�uD��}�{�u�^H�֖¹�G/�K:r�����
�p���UD�z�6חƅ�#슁�g�_׿B�ηb?��S��Z*�l��ic�h�@��'o����u�GI����O�X5�4˙@�{R�)���N(��@NqSƢ�ON�w�d\\�^��O����I�tqX
�^�.9��r��a��I��͌g)��@�%.Nɛ�B�����lfHέl��E4���~�}�k�cW�ueÒ�H���B���K��J{𠣱)s�a �#+�/Q�N?g=.@E���{V��ph��� �����}6��� ��������p�veٛ���ఄ7��`���)�\��J�'Y�����j��,ph�m��K�G�E���T�������c��N�m��J������aj��;0��D1J�[V߿+#Mq�2"�8JU�
8�NA��麍��Z՞��+e��1��f�Y����#~����ȷ�v��7�[������!��#�ŗ�f�������I��T.uv��"���	��]40���4w3%��M2J
a�2<���S�=O֕U�m>��d�������k7zH��},nv�W��r����o&��L��Ͻ|�c�M.�7�t�@wSs��Q�SF�O5��s���<5�xJ]��)�zD�B�r�ʡ�����}�UNM��u��V��e��wWS�m#�6T��T/���io&O�-��u�m2O*�pyy��n���	d����m�03�l�X��k�uo3ݔ��	����G蚜�-����΃��.hixc��QX����[ar�~����_�Ԧs���Q&��Ä���v�yt
G`C8�Y��	����(���J�#%۫��r#$j�WA�݂z!*��d�d�^�%$�i�l�z��Qz}<)�T?(�8Ӌ����2�C�X��|Z��xUf��6��z�O�/��u��$���PV�B�eE�Y���hP<��vW���/�&���N�!�����|T��p����0�E���'�be����%C��gM_"�cVP��	�8A�N��t\�:�
 3���S��O�n��ů�'�������Yi}!se�;,��8�6�(��Q[�hGtC�t��Gٵx	<?�;�O�S 8;"qs��:����2;f�S��1��ؼt��?1�@B�$	W��|;)ֶ��N@�`�ˉ�6����K��@�b�"�����d0���j��|��-I#��]�ȏ��Ϧ�D:;@	��ʊp�a��A��g��;��P��?��.{��8�o;b�����hъ�O*Ճw��e;�<,��[1�#ag�) g�>�4�9CHT�v?� -'�N��3v�����x���/�7x�G:�˄���������W�4.[�k´T��ݰ�fSr~��ݐFf�bW9�3#�p�V��e,6J�ft��h6qn\��Jv#�?�%2���ďӰ w���a��q#i��Z�D#������z�-�g��a���ExMeTu����)�s=�G�1qH;/�9"{9>	���OB�.��T�|T�S9���?��u�!��=Q����y�O	� H��F�e^���JS�	�sK��M[K��nc(�Y���Y8NAו�L%��{Hd��n�Q�U��,G?1�K���;��AB���G��2%�҉�l�rNmIC�Z���uJ�iG�C��Z��H�7���M��Y�B�e7~��d�C���6�ᑣ>+�ܻ��R݃<@�q�i�ߺϝY�r$���]� ��#�]�	�]����m�-�gWG~��ńj�Fh&�D�����f*l:�g�yÎ�.�� �7;@t��Y���[��bT�T���n��Q2�yU��&}#_��K�&wv�1�C��u��A�<�~��p�`���t"H ���Y@q0�So��ٵ[<
���;��4KT�4�s�a'����/''��3�X5�}��I�v���u ����:����E�$��ʑأ��<��+�`��za��i��p���ʮ�|;>vx�͎`\mɩ7��DN�Q��V!Q3�Q�:M;�:$���>sX���4�45�_T]�+�~��� 4R���Ᏼ�����xw����S~�P�L�	)uP2{ȴ�D��C��xL!Cp­��/��YY�d�
}o�F�9K�y8Ēn��9�]Id�>�N� ҥ$�_/�W���8��[M�^�X��?Q2��#��X��K)���X�i�8�d<4�X��7�*wFX��S�+����U^���W۰I]4��#rw\�#θ�#�f����-0�h�I��%��}�)/<Q͎ ���/�=���WaIgo�k��<^� l�B2���g�]��[�/�i���ڷ�3Di�J|���HAλ���Mv�؛�O��L�[r�}W�_��bg0��R�*E��E�qb[�%{x��B���ղ �Q��ز;�����	6���K�����;e�A_ٌX���U2�u�8�����I �0<�H0y7T��AbI>�OJ�L��Z���T
-ՕT9$��x���%V�e%F�6x��	�RJ����!�'����.����I���ѴF�R~�k�>77,�t��
P��D�^������:"\���,[�2��q9J ����0)e�ID�N��S�����R����^Z���+}w�������[�lǔ��/��k�u�t�� ~�<R0����J�$��9.0��nRE��l�xj�}��:�
�ċ���_ �JS6F���(�T���cJېv٥���dQh�P�L�$>nQv;=<��=��2�` ���vb�y�Uh�q{ SM�z���y|�`{�P�å�������j"y��'t~ �r ��^�����q%Ӵ�6�e��5W�Og%/ n���e�i)%�%�����d�q��,�K�R[��50�t=I"�@E��bp�xoM	�-Ry��"q%��L�� �c�<�eY�9��Y<Ve��X�xqR�����56M,� <�#ǯP��|'���ۿ*0C�bCʩ���$�%�@o������@
��0A��6�/�ya���g����΂o�Ѵ����FU�pW�f���j;tTG���}&�O)����/�]nƳ�N\�n�/Tw4U˹��x�UIq�{3{��S��А�Z�i��a��I�����V�����(�{kl�
�ާ����,�\��w?\uzBŦ��n��n,3v<c��U����m��><��2&l�ʵ�s � �u!Ok���~�>b�j�G_� )�}�7cf`��u\ü�x�́�$Ar|�Zd������n���i�;�V�	��p�C��'�1M��(R$ץ�"Lu�x�����-��Шq[���抬����B����
L��VrǨe����m��{d��Ê1z�w�e�H�@(�Id��?6���Jt�iQ�"��\bE��^b�C�d��9��3�a�{G��G�IA�dΔX������jug�1I��Xzd�k��Z�#`ĈV����,��	wp�`p/ͼ����,9}�Kq@���L�������H�хR?�T��$��}!�V6��>�������e�Đ���@GT���3�����7⎟l��2�^���Y�Ԟ�%���d�����t0�|�bE
��m�JUTi�<D�o:������9����)��K;x���@��hӝ��
�?��)����(�C�v�k�1_`�$�e8a/�(qz�ä��ظo���o�}Bp	m�F���L"��I)��<������"�W����$뇉��q)px��-B��\�֒vV���-Z��o�lE�]�y���'O�Qs���nD��R�Q�+2��w>r��;��#sCpw��������i��a���p`�*��%��X/�P�W>�LM�[O;�/h ���}�\;�it�8�����:�޳�OtPH�ݳ52���B.g'j�h�(���G�J�Į^"�8*�C��/�i�v=<�yW���� ���!Y��k[K:ǿ��c������#'}79�a@G�e����P�5����d�Mc#x�� S�M�+���&'O� ��t��A'@mH�"U����jH��w����m3����Tf�l�e:�$8oۛ�����K(�����WD�<VQT�\���4�㰡�W���x���IQ�"�1�����A�f2ޡi��L��#~���w�����4�F?��w�)L����q�Au��N�/L��[Q'�<U�q�/Sk1u�R�*���{�k@"C����m��)l;�س�w����DC����Iq���X�' ��	�
F9�)�Q,F])���vP�D��>�	��_�o�.8������iu�z�2���58ٴ
��KsF�]S�y�����\#Fͣn/���G��.�0��Օ�_����q�0����R�5�s��yJ>����M�^)h�Bm�3A��Qd�hh�@��$)���\J3���L��"b�tL��A+�ڃ�
UK�('�l�f',O(X�|�ۯrG���l�"#`
lG�J^Ĝ��(b�+��� �%����&j,�aY�X�;���h�h�N�	gw����U�$����hq��������&AR�Qd��b����m񖚫#�W�,��S��"	|�����~�|��M���d����Ȱ{�wϼ7�	�xw��(��&��Yi����/���)+N/��U����/���[� w����0/����Ů�NG���x�cP~��ADt��Ӭ�f(�#���L���d�T*Od��&�X��U	i��b���mV�=_<0,ȅ1�"�r�$ѐ��8Ely�5��5>;~������o� �fc�wz��7�0��u�\D�<�;�*�/�����G*�,.um�g��ہ.�p��O;�N[����.̼K��>���P��� m�o��.\��JV��2�b%hɃ�T�I�v,���>K�W���3~q<߻o� ��l���^��B�_������@)+\tdg�&qŋuZĤ3p�K�2�2sCJ�Ӻe����Թ�r���-�y'  �����}�;��|y�A�8y�]&gZ.�S���i��-�] ��Xn�S�\�堔������V$-l"�����@�L�%�,<� '�j��
v�L~�4��p����R}�<���ڢ�!����抩q�)�����)�ދ�-m8�r�Iz��;6�
�YJ]�A��)J�`O��*;��;- �@�t��/���Ӡ�ޗqrh����Q`��s��<�9�P�!�(�����F7��1��A�~��e}�!�$C�SD�6�����`�])��S,����E]������\�r9tk�S���i<�c����=G1�-Q#W3ýj�f4���)t[�sE����:&,:}��/D~��юP�m����s��Y�~ ���(��];�>;eҢq(�P���h�O�����F���A�F�`���1�X{~�!@���?Ԃ�z4V+n9"*}���1��B�^�����*�g����J�J
��в����t�g�P%"�
ӱ�ɍ�f�����14��s�;���i��K�����[�j�m��g~��&)\�Z�I�<(�rd"d�W�:)J��
v�ǩ��FzE��E�H�@��:c̦5��$d�&J:�<&D���wȰ	��\��1��_�<�LlB��Ŏ�WD/��C��\y,��^��Y�Հ��f��fxP:ك�(��O��q[�t�kqvP����Ż7�W�d)pb�%��0#����D	�J=E�/i�v/���}֭��Ѣ,�zL1˸������e���vr�b_ ���Ю�5�*��;d��{J�����۝�_3M��UA��g+����<+���q�� ��G�S��)��&ׯ����i�{�QIh�ײQ�����RU�> 2��N���S�8Y��r�'��(%�]Ҁ��Ex��e`�BU�A]�
8���ݒ6 ѡ:�R��h�L�L�<�Sb����4L�h�l�)6��Z���F·o��r���U��5u�"KG���J�3i��77%0�fY5��窐�5�"Nɩ
Zj����@�?���r	$�����}W�5%8�7��ԓ�~�]�I�`��	�Rk�ǃU�P.�o��>�ٰ��
����$�赋���zUKvv��I��o *��cBڎ��k9�1(���h��X�o"y���Z��9Dx�_�E2D`-Mc���%�B�{c&�N�s'��QG;�E�_�	�$���TD�0�߆��X~^j��8L`̤�:���C�ͪ��No9�� � �/%A��k°lF��E��T(V��C��
`���r�t_:ϫ��W�A�uL�V4/�7�m�Qj��ޡ�O+��ω�$>�y���ל�#���.,e����_��-+�u�[LT�1�O/�ax��/Ԗ�����,�&�m�;�k-.��R����?�)`��)��>"~4t��8ب��2�~��qv��1�b�y��g9_֮l�jD�s �f��7�A�A��) ��W�Xz=6�t�&xF[�߀��R�R��,%��|k
���z��!"d����H�9\F��]�3�/��L��y�����sgUT�1��-�ib�����*0�v������c���s���S�=��\�D\]H$$��Tq�r��x�?�h�<��{�<S	Vt�|�\U
��ioY�'d^�s�НZ'�6��]��{����1-�y,UԚ�ׁ�!���Тo�g������J����s~����x蠱�$$�?@�sYy�h�lϰ�d(�yOv���:����E�.�t���|���z��nBp���u����qq���׉�C��K҃0��:���O^(���`S���D������NL%Uy���C��R#؜�/���)�U�)@�m���7�,�溌��{=��/7C;�;]���i�)��Ur3*��;*C�EM"A�WF԰xj-F��%�T{�/!=�H{��4�o��"cx����.�O���,����f؉������z���W��U?�Fe�������T��˝�.�,@�`��Āl��M��qG�=y�5m!Ɓ��=���h���S��SR������G6�l�K����$�*��s��%(v�����p���눁E��ĳG2Adt#؞ͪCIp�}M��8���E�(�!��v?����r�����f���2�|�%�Խ#U�\1�A�a�1�v@C�W]ʂ�%#�/m�=l�ա��J:$W�%��L�uόg|iqSCx�Fk�h��be^Rq
p�Q� �t��Y�p;CҜ���F�_��^����s@_z�z�:��
ܑB>l�G�hݽ���Y����֬�Apڶ��uE��⽗�S�@�M�,DQ�$[�Qп��&4�u5<���@o��3ݵ�r͍bOD&�2%y8X '��x�o5:'�j�LV�g��39�@$M8J1��@U��\��7xa<������AI@����(y0� `5�	��u�C蓴Y&��xyL� Ff������	�hy膍��9����,څ�P UHO����H�H|uT:��V
f�`Kʷ9V)��K��&�2m?x�#2WX���,6/��C�ˎjG�Y�_8:tS�u؁�*4oWHl�^wH4�XȐx��6�.4��7���?̮�6\����d�m�.���bX_������%.{mLm������҂�k4������wb�7TBܢ�����ծ������K�y�[�С��w� %(�G�8_��ئv�Y�H�2OΣw{7x�B�j�)�P��&�Wg�<m�D�Z����u�`��m���9�Q�F�f>��}��ߘv�DM���V}��_K�b�/,���,�8��<,�pC��l�t�l�I(W1�%���r�U^d�G�\��|2�R\�����ԕ���[^��ZJ=G}k�JN#}���<��!A�twtL���x���=\�,tw^DFu�Y)c���Z�vrQm�-���Y0��X���1!N6�j-��%�,���3f�t�m�bG�G�T�ڣJ�OY�0�/Sɾ��p����nA�~S|�;��a"�'�G���h[��� ��;�Փd�������g���}w�`$������ ��b��Ceh���̗z;�;��	w����s���P�*���]����~�R�pY�D(U��)?[��5}�ɜ.��DƆs��*e[�7z�ݙVԟ���5�P�k��N���0_"!3B��I��C���qPR�
�D�s���0SaT����йp��<�e9�t>������4�,��O�?�[�)�tYҞ1�(�`z�V�H��<���m�`���e�˯N྇9SG��i�]\o��*��޴A�4�W�=�|���]�δ��~ۇQZ`�t��m�����,��Ĵl�䀩y��cSa3z�x�Ş�-�� ���������)��5�cn�i;Gk����^����?/�
*�2�9�DJ�S/{=�J�8����<A��.��)���I�\t�� ��TLXȜ�烚��'�Ϧ�imb	j�$�d�~��w���`Cw��J\�"h��ԟ��&"��݀��
���m��̋�!��/ϳ�*Ԅ]'�:�;�� �4ܼ0�L	v���u����Hę Ѓك|�����v� ���Jf���Sޟ����W7 �"�խ�5ohT^brT04BՋɥ�;CH�IV��F�O?C����`1!�'1�>����*i����V����-r8}a/�)`P]�	�*ӹ4n7�ς�xHc�pX��WV�����魚��L���x��Jc!�5xX���u�pq�ڭ���__%4��ݵ��#�s��Q��$��A�����8N����X�EvǕ�w�w��1$t@F��U�(n���ylGUܛ��)M�ojga~*�[�2���xc�w�����`j�0~�.�)o-yЍ#�p�mu��<7� Z�z�pZ�v폨rzN�_F���ڑ&�K�<A����I$�1~��x'>D÷W�?��m�vk�w�y��!�S:5~@�`�[ɗ�*�~�1C�RGaQ0�`5�{��8n6w��o�Y1�ڛ�ɶP�A�S�pƸtƍ���[�C�RU��y~��9(��8��&Ÿ�4,�I*xg�^bn����|j��~$-�<��x�D�(���D�{(xc�^wk춦��Z��[��_�镊���h
4�`I,�H>�l�|+aÂ��Ȳ��E1S�l�)�������^���������|�{,K{Z��1Xc�+�Z���ZtU���W��5Xxv'{�C����ɣ>qQ���^
r#�8��d܂
�g��(�u��~���Q�tg/�I9b��C��{P-��b�~��b9�������ܵ���l�cKU�|�ز������+�Rfn�*�z#���^L&�;P_�v����RZM�4K�*<�eYs}(���y(�v�AԬ��W�}��jjo/As��#�m��`*�y��%a�_i��<������?Z����s���F]��*O��W�S*H�{��L�Ϛ���U�zalpR��Y�"5�{��E���f%K������e�(�B��%�^��u�t�J�XU�3��֋�=����q�
�&Z��j�5�>��^tȏ�(��l'Ⱦw��e�YX�s�h��$@]�nڅ�}�3^��tN?�l��Q'���X��^� vԵ�~��+֧D���s1w�@��><8>%P�9v�Ѥ�.t#m�c�sZ����ɧ�c{��5?	���^d���,V�m�
1t2D�> �p7����qT�p��j:�R4h�a��v�~ƒ�3�M.��j9/���>R�M��O`�������0�6*M�p���W��7�?�V��É	�,uR�GZ��獬���c�V���?mZ�}�_^)������n)�|�([��S
������m�������(�����߇���#B�R)|�>��x�>�O�$/ ����>���M��C.�o�PvS>�#��ߢ��Yt�)��t���M�Ժ�?I�*��0���X��Le����i��;�Y�q�:e&rx̥Y\�Tv6B��Q4S�Tyw2�Y�%�%}̚V����jm������ZXP0�)HiRws�C~��8�>���Q'e~+���|@��7w����zy�Or��N("�t��O�1�ǮP�=��!�񓛐ס3��W�Y���n4.Hbs'�p��sˉ@n+�(��q4c��y�ّ�7�d�Ėmv�EM���� S���r���t:D��%�U��%i���ߛ뺴�X�.����>g	i�
#/�GU��o��ƶ^��6O�R ��!"���N��h6�_R��f�!��bfӒ�h3��-���m}R��q�޾�ZM���=�,��n�W��ܦ�ᑀ�(��`{ �w�A�H��:,���'�\1�y�Mm*�=YG2�eG�_�9�l��魹$|���a����w����C�Q��ҝ=��E\z�fֆR�ӑ��|n�CPaem�UXF7߆}nXC���/B	�j����|^�7��x�8��Лq���r��w���cĝ���JC�
��"���稾�y�`��[�L��rB04�Y�X*}��l"�e��:����H����!��ݜ�Q5�z܉
L�����`���]�����_C�6��d oT��cN��}���X二�Ѝ*�����_&������r`��PWV�����;����K��^L_9�6��3�0�빾̖Z�,;�S��8�,�x�����BO��$B�z��"n���**��f5RD��~�Ǚ�v�)7���ō�Q�(����9xas'�a
��r�]�j$��b	m��as���e��7XR�D��/=s�<�U�H��|�ʶZ�42Ҽ�Kj��ݝ�t�"!�؍UIG�@�NY�֛yx}��0ꋕ�25aeS�{���|����;7 �aiV ��K��eL��������}�dv�Ui$�]؟ bhf�0W��Y�mݸ}��}֖��4K7����L�Z�K�m;�� ?�r&�&��?��&�ϬBOZ�[MC��E_���탌�5�wX�FM�p��x�7U̻�/r��桲��T����d
M�A&`SB����H͒ۯ��7C�bL��e�� ��ծ�3�G31�H	&m^ю�4N�':d��P�w��ɋL<��� �>���Lɰ��T$�D���xr3 �*e�명_E���-R�3���Ő�8б�����ÇQ�^�5+�z���_Z� �(���YG�U=�7Y|T�@�V�h�Yi��F¼fʈ��.I�vj����<r�u:0|~����1c4�E)��G�� @�÷dG�s[@� %�}�r�&���L�H��I0Z�
]���U
S6�r[D�sG;�n�M����/�ud��x���[0^����嗑xC!4�2mu?����|"|�Äh<BpF�a��I���׋8�a�;`Oa�-���%\}ܖ0�ϯ�Ҡ�S�����j0d N����Pd[���?��4��)$O�$`�]�y����P�qۑ:��R��؃��Ʈ��w/����R�N�f�K3�Fu�}~���q.�U��N�ތ�G��
�s���օO�Υ3h,*��~�f����b���\빬��Ym!����%
�@/� g�	1*5�A�)HOˠP�Εy���~Ԟ`�$+����DVX�Eu�u���������ۓx�X����;lV�K̵�m�4{�K�AP�ag4	�p*g����'����;��C�B���|4�%��+���e�ϙ�T~��<^*V	�-l�
���[Em��\�f����=*�(^���S�N��_Y�s�Q|�X� U�q[�����Yna/ۗ@C4>H���?>��e�`w�s��z��y�>d�^(��*��J5�E�㞨lk����[�.�[o�hrk�s�K�7��st]�h��� qO�7�M��
[���%s�LЭx�[#0����->�߽�kUt@�p�'��<�s���:\���b+�p(�6�I����Io�`����D# �#���F��4���*Σ}��-Y�����T��I��n�M֋S�G�T��B.l���Nl�}�!��G��ZJv;ib��K'bU��J.�4Bʗm�� :E����;��A.��|��l�%��Ր�<<P����m�9�������l>�;�2�@4��4���i�wQ2gp\��
�n�2�	|��Rp��RV��2�\�*an�F�D�"U�S}��L����,8 ;�����ˣ|��9�V���c��lp�<!�ycI��j~ͺ���铽��8�� �Z�eJe�������� 3D�9vߐEj?Z���"4��K&g���sf���V�JG�1�*cD|t�<cFCr����x�5����Lx�W��2K+��-fe-0���X����7�3�|I���7���;����=���H��xa�Łp�~����@Ħ{?��$�k���x<�]��C|�����ߋ�Z�����8Ї���M�lXN���%
':��u6f����eF���FX���sMge�9��g����	M ��y�R�����&��S�a�k��ק#0sG�/`��e{���b��JN	������Վ9q��M2?�2X�NUx_2���΋���d��AKJ;�z�l2��!��'�U���AA�p��B�W]���HU��+��ޘ����I>��)����q`Qf�j�0,*��/{� �[��Ȗ�Z؂%=��V��qK�׫q�L�%���cݒ��F�H���@>Ǣ^��rٯ�2������Rh��.%Cx�C��Q��Zt��M�����w����ǲ�J`^�<f%�I���#�(|�Lѝ��( ��'l��RHTX���v��'c�i�nN�/���N,��ർ��+rD�(�m�g���[m�n�g׼�8���HU(��	R6�DR���{������fe���ƑG�JER�Z� Q�H�aq�v9�_F��jF��Ȃ*8�w��	ڜv՟��MH��i}����R�0���r&<�=:�S���\m���*G�Dz�͔�������S�0��B%)�w��NGƮ'4�T�sn��l�tvMzh����E,�)L��Dn���xm�J}�����Hs$��z�H�Y�_!����Qb����4�G�/�[�l�O!�/z���~��Z��BS�U�)�~DH�p(�!3�gg�ɉ��� N���r	0������
ɱ�h*�k�y��3�e���W,�J�ˮj��07�1�Ս�j)�Ӵ<��H���I���&�=��J�q���s���>N��ѯ�E��/3���$��E�6��S�����4�XJ����_��BV	���c�'�le0f1���a�F����.[H��E�	�Gʝh�:��ol$���1f�q�Lqu��o�}{1�/iɃ:�&i�k�DZԄI�q���/�O��-���,�B+�ӯ�_�8�q �-٘\�E�-0U�,�.�������-@�KV�aϯ	����]�١�*s5�M��y[s�yȐC����:Au�ѡ6#> Z�z�:�~_1�AJ��«c�_<8�|�m�C���ۀF�Uԣ&�$� �����}�ÍW���$��	�@Z����K�7�:���ӹJ�St�v�ƻa�?�Tz�,�aR�SNl��n̼~B���3'�s�2��x�vj���?���qj4���n�E��|�p6�|��P�_��Dh|h$M��Š�4NG�e�Xx9�$�詾"�͏�Er��l@���iusH&�&��%�;z�C�w�%s�~�4.�5�79aKfñ�i�V�8�|C��c��2�)f��}��'H���N���>�-RiB����P��>�H�O�/'��V������e�qF�9@�&�����e*O�JkgZ�̢
er��M���@�Q�3/�����x~��%����?T�6�j<<q�7��{?jȂ�T+�9��/�6�\���p���N@�Nb	;|#�JI�;q����Tn��S�"Ѓ,ƥ
A��wB�ub��!�:��/i��(֓�m!�4�J��������L�kk��~����q�1�/�),��<��	�������[H���I���ׯ~������A�W�˛#���E+q
���F�/���0YMdtq�Ng�2Uf���Z����� <��a�v���µ�IX�Zڅ(�,\E!��A^�@
���yc�X��D��¹V�%�O�/r��]	e��{JPr�,�.y��ѵ��A�^�0�E������Q��p��yGz&G�h��[ #�Q])��^r���V��(W��Y�hNvrF'tIN&�1,e�\}2,AE׏�P�0k���F���;��20��JNg�H�n��1��w£�#��
3'��'�l��ځ2�~.+�=d�R4��44I:��pd��Џ��R>��&t�Z+Xo*�� F��S1�����/)�It��&�.�`���Xk�ev�7;J͍ym��: �6�/���-���T:ll�� <
gk��5���Z��(|�U�$��ؿtd��v�EP�f��M��D��o�T��⣖T�����ߎ]Dŏ��>��L��Jz62�J��lp�P��AQû��u��9`^��f1�T�,gz��k����nv���������5�Di�soc���%e끇;�/:Gq��,V���j�����_2	��'�d社�CIBlے��ZgZZ��Łخ��$?�S�&U�eY�\b?)e��۪��Q-��u?��u��c^B���V��ԴF��A�BQ*fa������й�1	i�o��㊆���,���Rr7��L+��q�q;��b{�*�Џ���YG�ݵ|ン@�i����vM��'�*���&/ɳ�����JCe5=��s�����s��L>���V�P���	q7�#�ݶ�'��������b,�������n����g�g	Z���Hj�M�]�z� �	�I���U��]6�Xj�W[��y�l;����,��}��w�Ü���}�#e��[p�OۃZ��Vf��~ ��(Te����~�Pi��G���B�\���}V=�ʿ�0��0a��F�a9�_S�/lua�,�/�qZk���d����!�DC�~{?`�V�J&hF�#�D���L�w�|�5�M{�x�R�xfbs�H]d;s�imX��E_i=�����Lx�x��������c��??E��>�zq��sk���0!Zqvy��r(D+�?i*[pk'c�r�k#�(�C�7����ro�t)�b�pAD�8�+��/��j��
�^'Ef�B�e#s�?�ܥ#��7�k�n[-�,�hB4�}P�d��T�ʟ���%�`+�1p)������݊v����Hi��~�g�C"N3wM��ޕ[��OI	���a����+Ǌ�}�y@&]�E�c= Q�oy
���l��#��据��p<��Xf�49��ݤJ�˞�Z�1;��웝��}���YrG�跖.R�!�.ѺF�6fu�� :�E��|Yu�����R����r�b��x��� Ep@����Ը�t<x�������5��.��<�0���@Cr-��m�m\*���`�v�?�Q�� �1#W�H�_��K��$G���=�,ʓ��c�(C6���$�ni�Z������iRN 	���}��Hu���|�I����F�*�`gS��bS4k���7m�����3L!A����IE�&HW	��e���&���f=TAN�P[䌝E(�#��҈��Z�Xb���W�T)I�|;�����]��� �Bˬ�|���p���?���D4�	�K�{�������SN���Oͷ�Ċ�J>�w�d,{怳�T�{ԮQ���t=�O�Y�_3�ْ<��e�Ϊ&�\/A��5�ꅣ��TY�J-G\�	p�̊f�YU� ��X ;b0�_|~���Zk7�;�c��������l|�:������b��+�)6|�Ho��U�p��Wq��N���yM/�x?)��`*����t��97VJ�����<g�Y�V��|����L�E���I����'���W��f����&r�o;]��P�h�pR������xT[�==kxN��6btK	�-4/x��|���,k�Ӫ�Ȯ ?�BَM�F�m��_�O�Ao���6�F��y��l�7?>��:FYÚ2��@-fv�"��7%�!"�����)��ڗ���rV90i�>�W7|$Լ��ب�ȥJ/N���^����)F�P�����Θ�Oc~Տ>{����'饘�Oo�f/4%W,O�S����;f��@�I��?�Vvp(�Zp�	�"R�'đ��
A$���я"��'���3���$��s�Q�'e���;e��+B���܆!uEv���u|/ڣ�01��;�H$�}ڻ��X	 �
.K��7Ɛ��=e�h��^���r$鯡/��c2Y�t'v)��Q�I98>U0�2��H�v)1�	�;-h�C�D����܏ǁ�iǢ �kM����<[�Y�?��m���V9��=���Ķ�5Z���w�A����������P�_�/�`G?UP<�[���ъ�h�WG��F�zYЍٔ!Y��^�Etf	��s�Q`�<�M"�X������������<�36�� ��֞�w<���҄�|�_	rZ��P���jr��O�R\�r$�Ua��y��v�M��y+n�p��y��H�LVe�R(n����{il+�k̽T�H��ք���9sN�:��Ҵ�%_e�)}�s_o��vL2�$�/�x��&=<$瀧o��u~��/�eC�!J��{݋�����������h�8����VG1v:c<�Y\���Y;8:d�-�=_��`��s��~�@��)p�H�ā�q����5����C�*lr11��<J�L/���pT	��S] %\c����3:7>�(�D$�@����W���`Ȫ`/bz�ȢT�Zι.�LV�K�p���	�I�:��4a��u��lF�bר~�EX�)��Y������"��\�!�lB���JҠ��gz�@3�ߋ�X�\����J�Ə3�O 3J��i1*��q�����,���������	w�RhM7���D��n9�pJ�Owh�Z���	u���i��T�p�F����m���/����S�_Ja-��xp�KI<�}M�L^!��F�	���:w�O�D\����Oz�&�A��T��Aw��M�����J��S��A��|d�D7]Ь]�<�/�S��_�{��5+]��Ӭ"%jj�<��%V�v��'�۟��F��I2C�Rm�����<���f:%C"�� �9��KE���NMf|6�|�Z���6��n��} ��
��=�eo���W۟j[�;���uy�W398p;RD"��ÄxC8-z��9W�{��=x��Q��}�X�ց�)��V���'{Il��vM���$�@�\��'��q��D�_jr=Ƈe_Hώ��J�g�Q ^zJ�����ڋx1q��]8���,n���/v ��\�o�X CR�J5!��<��]�&V�L�i�(���ڄ�������`���Z�ɱYTo=8#+��߽�piQ�T�b��|c�W>e��X�'�K�<ER� ��tR�w!j?�C9'H��ɷq�����?�n�6!{pι\���XHvF�1ȕC޾T��.��$�2	tќ{M(ԑ0�hnh�D���@A��h;)ʳ|W����zؗآY�wĉ*�Æ��1���#�=C��+~�K�z1�mCgȚ�atj�ѫ�j�\�?�#Ҿ�q����E�?��J�����=�9I������0i����z��9e�=lG�Y[���|8z�k�E�c'q�1�#7��Ú��N��Z��P�n�x���r�1�y�i<��5T����!�F��"{=Ac�f�!a��^�1������^tQ)�L�,��dJ�Z���Bn�@ H҆�0��ݜ�až�J�MmWF�;��;���Hh���2t0t�W7m�":Uj�	`���a���1] ��.0k�:P^��V�������+�����e�M��7b�!��!�gx@m �Q��^<�a=E�
EU��
hǛ*
c6�=����@���B�f�AW���0��Z��v�@�5�G�#�V����E�^��z��u�n� �$�H���on�x���G���+�!�����`K��~��SV�1����'�$�)fF��L��#���{R��'�H�k}�|a�����u�ĉ7洃��`غ�W���`����Ս2����;&�Eb���ĤQ�<��8I���9Oon�T-I �; �q�
���ƚ��hR�}��?�& �6�>Le�x|E�O�l����Κ��5Et��x�a�n�&'f�==3v"�h �Xw��}�_���6��y�z���� ��i_��ȣ�� Y�)�N���V�����!�
hN9����*��Ee�N���K_�\X����fR����C�;j.S��Y:�oI���9@�ʡ$�~3�R�.��Ȱ��WS$ G-�#k��'7|���1AeX�7h����D�º�w���W[����m�"�VZ[ݿ�x��U`��(���9���"�\=׊#5s�|huee�L�$T{l���ۺ���	As$r²����v|0;\	�k�&C���[3����}g�耊����ȡ}7��L��	x'J{0a�ގ`ӿ֝�Х�t�L<f���]Fld�~&�¯����nb偸�Q�;���I+����2[�:�!4�xnp�NB�ѡ�,xe���T�-c¥�붌c��X?�W�0��;).�2KmO>�@�ZPN�~�y2|쥗Gڪ�8�A�ǀjJ��c��~F$�g�:P�[�ڃ	��U�<R�I���k�!댲!پ(d|�VX�fU^���9b�ٕ��	@�O��J:I������
kF&�Oיʲ�m'0a�>%D!���#@!�R��� ��vy{a��b�'B���a��a���ᓕ��,��;Z���e�p��K�$1pu�×�R�'B�F�H��K��Z"���9�p�i�]���h���W=+����[������-Yd�R��J�=?o�u�XJ�Eyy�� عD�X�g5�m�7�`!�~U�=�:g���v7�-�G�����Fr�B������Jf�Jw�c>�9-����$���nߗ�[\�A�hu��*��f�6g^jAS���7@-�Dv#!H���}3�)�m��ڢ~s���-�Bc_�z�C�y�3J����p�� �av�J�NQo����$я�ذ����W�����M�R�P���F<=A�?A�z�!ڽ�na	/��M��G������F��G�,0���Ģ.��
��pt�Pgm�L�L�#���7�*���9���r�G�7­�_;Z��=T���=���t���-� ]PyUM
��AW�bYȲ�/--�N�p�E��X��H�,C�l"�C�������7�I��b8а���<�<?�ӚԾ]��체K,3�Ũ0��d>�{�����s�c�#�.׼��9i"
�@N��6�!
�I��se"��	/��v�U(/���D3�.$Ѐ9 ŭ9d*���Q���Sm����q�A!���6,v�K�}$Eˣ�.�|��8|��r�K�� 2��u������]f66�W�ݚ1�j=���E�[)3�0ϠB���<Ja@�.�c�kZS�����,��?2]S���X��'����	&�`.�i����G�#]�B<8~�P��뽗��Z�,�����C�w�{��|����� ���S:���T"Y=��>�)U��B�����_'Hv�ؠ����Z�A���E+�,������`RZ��&!)�# 5��.���i*.�\���3�^q�}���n	�5�j��o�M|��2�t1c@���g;��}��^R+���?��CUS�U��0l���>U��(��h�`�tYu�[X�ӧ�)i �V����<��@�zfG7Rֱعs*�P���3�ΰ�棳1�1W�B���F���u�y$��D����`�����^~��K�$|�.�x{/�C��ؒ��ڦ4^%Y���� C�M�Hj�����_/;�w�� ��yn�KHԸ��(�K����&;$�)d��P�(Z�25�]��w�z�GD�j|��'�ڐm�$c)��g��6&�ƨX�����ߚ*�Y2P�����k��3"Fk)�[�v8��"6_���!Ӡ&5�c
򠕃H���.=�O��lo'�"r_h��S��I���/��!
(Ö��:�HZ��.rW�
�j��\�����~�hP���v�Z�4~�)O��׊���Җ��5�;��
WUҐup	M\Ӭ�5]�XJ,�O�;�� ���_��H��)��E���>�:Ef�c��=�Q���a���%Ö�U�3�����>�\^'U�)
����D�_��,D�J	�E`���� ��o ]��]"��_��_�Z%���:�mO�ӘKc���^w��-�܎�4�!׭�'�Ҝ"�Sk�]�nE=�YѤ{-�Ie�=����|���(����K�b��g����V���R�	��v����mS�}^-�d\~��Fq7��
�%��;��3 I��?�:�^=�U�5Lt�k��v<�.��u��  ��JPRSƺ@.p�p��Agd#����?O#2��R�5�dT�'�"��Z`ȸK�� �q| �7zu2O���IJφ�+ImV�I$�IGJ����p�3������T6�����(�q��<b"��!�����m�龸/��$��m������-.UvZ��8�'�Y�k��2ePX�U�?2���i��a���7.���+A�#S	���Q���/ˈ�AO�.�<����Ӛ��ݣz�h��*��XB�cL����.�c�@�
�廬Q�">r3,9A@�O�12:%ܬ�AjN{��;<Q"���u*�y��{�:�(�����;���"�'iʎ^i���)q�h����$Pc�%5���Z�TM*m�؏ƛ��Ēo�:ǃy2}j8����!��g�8N�����kĪ���1"�x���o�x}1lD����ي60�MJS?�R�QF��I�-OU�>H��q�R;��o����;ܩ�J���q\4�[6�ü�A˼P��8=Jg�{�N]e ��Z��r#o���ED8J��.���v�hͿi�&���O�,(!�GL���A�v ���C��V�9��c�R�r��?ϵ�C��Z���O戨�<�?8i@�S����6��w���s�h���Ln(o_��;�$���?���.��38�}�oӐ����yr�K��h�N"�Φ�v$p��2�ok3��@�!!/ׅ�R*���9�t�����ӹb�+R�e-:��qMg����r�>�#a���u��I!�>���Z4'�
Ǖ�?8�5P� �F��mP,ɒ�
q,�H�u9��(�_7K�՘[�`^+e)z�bz�)����+�U��يC�ݰGp��6�z�~��g��:��D��̐����<��(�\���xT���!j�=�#��^���p��BEbS�0T��\�� �Rr�*b����u�K�^l�gt?�yp���1aG���eY>}� ���+=���^m^���O�\�\�0������m8_�U\�k`�[;&�=��H7~ƎPr��6,g��W����d��&��^s���,�;ph"}o^�Ӕ�q_�G]��g�7Ϗ8@�T�	�|�x\�������~�v����t#B F��R�\fkG(EU�+H1������y�������dڼS'<
�b�[4�>3�b�&\:s-���Q����Z��H�4����غ	��^��k2�7w� �s�������d�D�����l�ѵ�:���4�a���rn�������o���XDU��r� �i%C�ţ�fa�B�M��<�}�Nɞ�Ҽ]5�A��s�w���5E��N�̗��9X,�\蟑�	�[�B�����XC��$uy�Yʍe�y��P{�p�p���H������_ɟ68��U�a�8eL���h�°qON��Oڳ�u΢�C�Q����^~��l��uoH�@��;*��W��p@����4w\��J�MB��b��/uI��n��K��;�͆;� ���%�Īy'C�˛ �9�vvxX��0����ۚ�ȍbцB{[+j�09�7�s<�`E��HQ�U��0�yz�s���v��N���N����<����^R1{��ˢ������:@�>�p��s�	�1�;ߒ�ݠ)@t?�� P�s�Gg�h��]l�_5�50٠��9�+��ض\IA#�bOޒ���י�$�&���k�Y+LI`�Z�7�����oN>[cq�$0����TI�c���@s��"�&n��ƻZ�P.��2Xj��ϭ�u�~Z3�"��e����W����-Bۚ��y�rHBc�%:�Gb�ݑ�~�f���?��mUw4��U�D��L���&�G:�e !Ե�̐b�J�k|�c4S����3y�d�?�Y�3�eE��kXV�Aϗ�4�;6$4Œ�K�̔�dq�X��q�&��&o��q�q?F�lle�Q����&��e9�R�Q'�nF����ϱ���֎ڻ��M�\|
�GI�y�EQ�$�V+A�&�IΔeo5]���ߊ1��Wu	��h4L�i��k 	$z�)!_ho��jⵃ��=8�MN�Cx̂��@��z��6�\XG\O���bV�0�P�$�UT�yٺn@��Ƭ+��u�bj�5,�{�G������0���78^Z��z����L�*�7�Lyo�!Q3��6a����o��ع$sg�#��r��uR~�Ê!�/T�ջD��0(� Hu����;C�[o޵��	g6���,�v���?ub��-��1��*��7)�3�(�E�1���{G��z����Sɭ��)�K'��
��8�������<���x����T��E˙�g
)�/#����c�����0���%o�ĎC<�1I_x �#�sb}�p�&#�hRȤ���@�[k�>�L��������� [Ah+׼i`o3ag�w�����Y'�?y.N���D�3_��#���XD �sO:(W�c�ڎ���`�됮�lFS.4�����A.�\��6%uJ۞����aL5���}�����J�r�ף�2���^C�Qzn�]Ա�ɬ����O�L]��W�lޅ���,K�)G+�K����zғ膺bo��ӔG��Ӄn�p6�a�$�����"��S#KVb����7!��#r�i;0P�[�ߟ;�3�}\��w��f�o���}�q�T�8�ۇ]�l���jI���F��
�i�	Ao��q�	B"��={����>�B����lTI�C@~��/�K�0SM�����3�A�"YvbpR��=�8�s��Q��J`G<L��dh���4��M:J���$;�M<_T�����V~�658�k��<����N�&>�i��.2Lr��p�tbNsF������}vw*7�s�'"S�:�+F�ݠ�WN+�T���-;�9C�?	YЍ+��knf��=�v�(��@ƴ�:�Б�Ms�]�%� N��Rd�	mzWw�c��ҫ4 A�1�ftLRUܰ�����;�%�wz.sġ�tr?a�y�?�k=aiZ�7����K!�>M�� (h�t��61�BX�������_����ǁ�& X](����BRTW�S�?�8Í��j}낣�>NI����؏�S,'�h���v�E�E��F�Y�`��S�o:c�D��%[�eA��ʏ����]@2�˜ � g�b�B���x�)a��8̃E�8�L�lݷ�{��o�g�=,��+��<�}� g!�����W�p��
�nE��qh�d���|.Ҳm��UH��F]�Rmnr�����	 K��cC'L���V��+�;������h�3R�a���eT�i�6!Ũ&K����m���m��d7{���	.��gBcP&/�m��ΧUo��P�O���x	��r�V�I��E���{y"ye��R�wB�;�����q;�:j'��Gl�-H�'������9x�
p�⢙+ƋPs�fc�-x3�Ä���Q��ЃYfF��ݩ��]�حmM��	�9
c���S+�jO̢�z�)�q�V?R�]�-� ��2F�F�����}lC�a��F�u�u�����'qU=d��L<���T�V{����(���<}�Yn�zB����:K���B��U������v��z���v��>)�+�,��l#��D0�q��@9$'� _���Ι��x1< �y����$��u�&��%s��?�"�$a�D�p�Os��<����4�B�{ıi���C���7�Oz�@�<-��Ў���_A��ʹ���1{�o�I"��a�rKp����5�u�v�`J����)��XZ!C$�[��#�1��1����{:t�x��/���K�TL?S�e�$�ɧv�~�� {���_�(`z�~��f/�>�ݮh��8Og�^��<0+�M�A�������ya�`��� @d�:�xl$p¦��\��(��� fG�����х�!��2E����
Y�3���v����Њ��n�d62j���RL���_���V��f�]�"G�T��;f��A��*e>���>�'C��k��9��oM�Q�%�:�W�� �@_~��Gg�1��L��{�X?Lw�u�P$2��W�V��I섒,đ=������l�c;��w���H!��y�gOF�4�a���wh�tҡ9P�O���4�$>7;ԉ;�ZREEҽ���yE�^�.��^ĐY��ؓ�=�e�t�����[���Xl%u�p1si��#����k5z�Ȉ��5f|����-QCw�[B`������9^�T�
c���}-z��&�ߵ[�HH:��_/�ԆK�QnPkM>�[LS�	��!����h;%=N>����>i����ǽ�*��}�W��ݑ�aD�-+	V�&��̠�>zω�;4n�SH��(�ї �1�k`+|��g�Uy�9�e�q�N�.��7B�x�"�D� 1	ҕO�;T��	^3as,�����;����#��
-KM�C}�6�/E쌙�\JՊr�}?%�<A���"
:?���دK�|=���̺b0�� �M�7ȫt�t8U
�<�B�q���i��*kXf�M�s�|����[�~7��#��^�QB�q���?���Z|>h��0���ٮ��O�5B��AI��qC��1������T��̵U����fJ��j�:��l�,g땗��P�!ڟ�lp�@jv���X�$��/y��}�xH����M�)G��Ga�A*<�+)0�xe_�_~D�)�HG0�׸�u�P�k�0+����3��R�!n>W��*h��.��gB�)c! -��>��cI=�9w�./�	/-vZ2����׆�¯�|.�Dٳ~�H���7��=����0��g��!�[K^R�o$M�!��*�������?e���pqpw.Q�4;�E
�;/��$�|�D<��CkQ�q!G3Z%�Y�P?C�߃Քk5�`
��� @�5W������&i�E*���.����:{�tk��WCG�P3ʯu�����0�'��BHZa>w�[��[�:��,K�ȑj?�5�[�����:��Q=
�,��L������[���q�>�^px���q?���ms�N,&"��g���6���^=���u"��kC�Ca�޹��u��;���F�'y����m���x'�w\sv	��p˾9�EFࠑ��u����M0?��H�l�C�X 2-q��a!�-Ͷ��ވ9&��,�R�&:�	kr-�[dx���wbX��z��,U�qrj�7���q�6]֓�<���]QA��(Tj�n%u���P����2 ڰ���ȇ_�	�����U;E7o�X<�_Ј5| �"�pG2���8_���|�h�0�%��V�`V����EWd����{��V3����K���#��� ���r��y�{��{^��S���#:;�����aR��Ѷ���e�f�V����=���-vC����Fx�m�p�}�ޘ9�-������XMR ����^���ѭ�g�pb�-����D��&�j���оceA.�թ�S�L���p`���O���H}#�	$F~��+=���QEGfAq��n�WX'�h��J�M<����A��ͫ�������s*_�%����sY�;	�΂B��O%#�%��iܟ���t���u1g��8�<�5�r�����O���2��m�˘�
���k�2�@��"W��W*�e2�Lf�y�FV5Rmk��7h�)Ev_������*l�L���l<��{6�����M���IP(�tIkD	�IQ��,���z�+���JH~��W��ﮜՁ�3<v3U -:��  l�������)�� ���2����n�Mf���jL�g��>a�����1�+���տ�r� ��x�3B?!��Hvb+��)�Rm�M�z�i����^#�nqDx��4v��{`�9��j �����1�T4AL��DnԑJ�|�{tZ��j����y�O����)�F[ݾ�������}���iU���b�`y���� %`P�^��� G���s���j�{�&7a����g�o*d+�zNx��P�I_K
���0�[���^�]��n��-������;Ć��g�T!4<�E���X�+�>�e4CH_T?��G�	h��(%���iTe���|��i�5,d@�yΡ�
������u
��i{���Ѹ�%��e��%UP�sA����Ң~�?_�������(?Ӛ#��4<F���b�$���ؖ6\r��ѥ�VNc�N)�B�OY�"�w�'�����L��Ν���2U:jR�_���.s��s6��[�tk��e'��\�)���f�j�?�|�ڡ�����{��Tq����6"Lނ�W9���RA֦#�ڀ��?=�*���?]��T��e��M0��"��� i0�ziW�t�~j�W�.�o�^������Ƙ�|c�,��Lhx'�hv�����x�{m���V�
P`߼��W��A�U-n�c��S�M,�%J
��MR)2�zT~'E� ��8�7=�a�f~�&˳�>����0������۵j��B;�-�t�A� }��!��p����'�rM���B+0-l��|Qw,�Oƥ#b��!�K�'�*nǤ-���J���0S)���=Du���1�K����{�5٦��u�>�-��W��֌��&P9����M�vʌ��t���5�>�t��6оdy�g����9�2��,]��QHD�d�asX/2������.�O���g���o>�5�9
�&C��k9���ζ[0/9=� �]�p�o|�<�Q��{�
|)�
���&~8mT���F�vߟ��6�ȓ��K���?���k",n�I�a�Ԑ_#Tm��y:������U3�#+K�G[��7�3�Y��yBԿ����h���T!]&�s��6�Ȏ�#�Ar{�7P��	�?�s�h5��N+���WMY�}�m�M��p�����c;��e/PX'�G����Y���:�WI�#�Mcƨ��2썐����=}�@���60��n``K'����ML	B����OU$9ϱ;��;���k�b�Q�<I4-��9Ltkd]��цoC�Z"��?gYc���z�ei\w��z�=���c+�G�� �_�Ά�a��6����+���P3EE�#����(��{ ;1�>P�W���&�`�u|
@ZK^!qjv\��M�|E�&��e�Y%�0s��!�w�U�o���bzw$��txU)�'�	6��w&�,,H��:��os-�vC�@VHD�9U�֘���X�F?צ���lh�C����2��S]��v٨s���m1,.� $��^���@[u�M��������r?aCзmC��Y��[�C
���-O�W���ǲ�G�6���ar�x�iۻ��J�0����v�0��5w�h��M}>.�K����2F7wR����0�Eg_��h�K����Ƀ��foY$���aԱt�)�L���Mh�f�}E�:I+6��8=�dsG,N�T�s���U��Eb� 4Ş,y������Ѳ��oϩtE�r^��T�����㡪�z8[t쇠��>2[�ֹ4�ԅ��ͺ�����Gu��
�VX��	���7	�:��(�M�&.�����փv����`;�X��Q����'���}"� ?,�������)��1��1w�f�^�!4���)6��`e��O�N �u�q��{�㎋ �CK����vo�y��z�_Rf��*�2�̄���8�k�0�͹��4aOX���I�y�D������(U;̯A���������g~@,�+~�I�X���X�*S�J-���5U���-δ����'�4;IvXA#�o:�ǌ�S_�y��LB�5 �0kH�.�(?����=����=�1+1D<ϙ=W���jD>��B�p���ܢ4�Q�I��ܾoLΗvok�E@`�&�Lv��/�?����}��^���ʄfEG���$)��=�0��6�����k)2Xq�D��'Ԧ_�-.n_Yl�	��߂s���iN�0|�)����r�mfy���w5�˾����d�^���j�􃔬���۴����{�y5(�-�Aj#���z0�1s6�4���6Ĳj�%E;�ցD��8��{P����:�?�\`��!j��gP�2�`S�J]Zѝw���'�Lq�6F�e�Z0��ST���s�#�l��5N�<��sc�9?ǒ]H�?�!U�<��e��a$�b�{���ht�~O��SoنE��i!l+�ް��
�7�^�'%�g?ŏ��+���k�2B��%T�z�s?���u1ΰ���߭�����zˁ�����Ju4�7`�=J�i�M���^@[����i��>�P��݆$?��%�z�(&��N�!�_�<��Mz��	�"����\�%�I���wa�����7>t,���|�nwz�K��2��tV/����YV��g��YD\�[����v�6�`���z�)��hua�\%7��g�cB��,�z��43�#�9��9�*�n�Ba�K� Pb�������D��c\���(���\$(�B&�u4-�����Ƨn�t�~�*��87�͖��Wx��mvR�X��o�7,Ľ	� 1��mv�#Ip���O$�M���V�ś3��j���az�dؽb��"��P��)����6��J��YO`�������*Og#�;
�=��R���{����aV��D�!%;��SoX��5��o��ԧ~���n2��dP���d���Ȧ�����x3l�B�Q71�΄��>���NWEYc�rϛ�ُ<�;�ʨ�}&T)�Wi{��8g���K��[X�>�߾më>�^#��.��n]����eQ������:z��P��t%���<�τ릺Y��K����i� J���x{F���٫�'p�.��C�tlf!0�v,w������5Pu3
�mO:L�sL�H/wf��]7�[:u:7.X�xC�认�vV=(n��X�y:Xu;"���Kw؂F���$[��D���� ��m6~#�{���&���rZ�+� P��n�<t1��7�AG�f�,�1����Ù�be0�<w��Ҧ�s��y�s�=�p��܆]�ơ��xa��{�L�~������#"X���a4�%�
��o/k��Pp��ŌE�����f��.-�)�*ry�;|V=�r��gm`s|�(P��Ğ_!�ȫ�dB�5%��v9��V�1�&բRy���]�fSq2��)e&�NK ג5��F�K�Twdߋ��Li�v4+��	�'�ڈ1_H��tIN��z���W~N�;��>��X�ʜ�<�l��Rm�h�-o������u5{x5���F�����ީ�<��jD(�&��ы��[�0�%c���V��Z�\�:��T�%P�yx�������(P��M���W����Z����a�K��B��f0�vw:���Q�p�&dTVG_5����X@�H*�X
�]@�_'�,R��,�S�AB̰BtەU���y;��ʸ"�yt�����RND��i�Z9����K�֭�n��E���[o� ;Z6u0��ɠ��{������Hw�Z��N�3��7>*}_�D�F�tW�
dG�6&{5
���ss0�7��i�j�~����.��L}>+{!/A�'�3N;iKZI�����G����f�	��-�eDs�/���L?QY���¥�/��,5��Ө�����?/���a\C��A�Y8GVLfu��!R���(�z��'EM�u�?v�ʀ�>V�7�D�u��jcc��b��Ln�̀���R|��0���<��WW���Q��Ug"l%���9Vd��h",���n&��h;1K��t�-�[H\����.kt�R����������wH{�)%�����������*�&Y!<�����m��M����_KH�
7,A�\Q#Di�3�'XX�JkSg�g���T��������u:E>_j��X/�5Q�H������8;uJ����|��c�K\1����v�b���A���fΊK��3��記�و0k��,G�69�?s{?"�I�+է��.:D]j��=w���,��LZ!k{��IȈ&��H,�A�bP�JP��,ZӖ�������!O�:�P2�h�x��%�Ҍ,C�[�8��#�
�ɱ���;+���u	���Ťĝ[�tKS�گ���_�ױW'ܻ��#��M���)�m^����ٸ��>-L���	���G�H��x#�
������5DP�,�p�r����� �u[�|��R�.�/��R{nS��W{���1���,%;�evO����T����<��yА�G�� ���2��N�w�s�Xm\�xJ�@�[�x�Iٴn�EeDĭT�-�ǁK���J�3��?J�<g���$Z����&���}S�j'!���<�A�,4[|c��3�ݬu������u���W�u�Y�Q\K
�� ��6���=�.n�!D�/���Z]�K�Tv��A�6P0�$�ӄ����畢�S&C��U5�� ��XW���jxdUB�rW���o�mK:��YV)�8�$r�I��8�����m�Q�?Y�����]}K�d=+��+&w�q9W�qV��Mw�1�h�=�a������H#���_�\���ƈ��ħ�{;��5	��8e��;(����j�g_kA�$	_g{a-9��"-��	���2QJq��^��j��A��-�6MvZ�+�y6N��N��ފ��  ���Lo]]���* �T�;K�.Dr7ϱ2�&ɰ�P� 8nq�%X�鶫U��~у"�Koe��6H��5��W���H;���L-lr�]�-g��	L>�ײd8�'S�q[qj��DXװ�f������X�S�v�~{<�T�ͧ`�p@DČ�B}s�N�G弍�f��`��mq�8�#�(�ۅ�Vj9	��� 1f��͡5@X��*n� ~�+��@P'��$��&IiZA���Y�b�D�I��όw3���B~.:���l"��:ڍ$On7�6�|G��ޅK�[�˵8�)-ք��d��ٵ�}@���MD�s||�	̍���� DH�^���a���w��.�`�xg+`ӵ!�}��P�R�P������D�Ên�湮#�)�+�YL�5"�����-�������"R��R=��D���O����jX�o�
1�c�&>� ��1�R%�s��_��!��>-/����Qd�9Vˤ�ǆ0%yR�&Ł� }XFB.�f��|�W#�!;0e2��	x5���;������p�G
���V��ѵ���,b!ʋz�4�CRLۧ"�yD�@���i�<�Q�e�f�r�/!�P�&`;�"(�W
X�Ƥ�+Ґ��l������K�'aȓw�~
��Z�~��<���44FN-t̰<H��|Iw6�l���m������njK;��N�|k�ayd.a��g�GU�f9�	@숚Dg�Z�Θ�>�)���$Ȝ�e�>�L��	,-��x��:�����l/�U^�79�^,U��t<J�@�d2�M�c6R��V�%a�LiI��o�7��k�a��{��W<Ҁ
���Bg�����e)ؿ�.b���吶	d�a)��٦�ߋ���u�n��Q�1�[:���6��JVXe�܆VQ��K�1�"�$�Y-�����E�*����Y�(�+Y6�M��9��������t��⒌�a���NX:������Y�.��<�k�t����q�0��A��n	~P(�bk��Ľ.�����P-c���Fl%����o�ߝ���M���5�4�jY��(��1��N@��^��] �mH�~8=�{�E�q�X&�k9'�M6�7E5�����^>
��~6�{�X��*�3ll�oQ_gQ��FV�N.�k�w	�������~���i���A��A�mP��&l��@^b���Q,���e��T��o�C��ɶy�N����EL���ث�45���I�RE>��-"�]�vMa� Y��`�y���r��j{k�*`Δz[xxo"�ƽƧA&)�o�P�蜘��]O��U"&G�׽@8�\�7'_(m>T�a�ϕ���>�M�p��ᙏ�{�e��n|�/�1&6��+'"M���uI��y	��xa��۾���-?�L0U��)�֦�+��*���^��Ů�q.�rA�p�3`����@ts�4��F��5I�V�X�N�a��IP�Q��x�Y1����E���82qK�Z:z���=D���0�9>5�{��	�	k�}Y"�\��[�:!��(w�cf��?��6EA�HF��A�<�]���F ��\6È��VƦ<�*�&�JZ2�	(��Kh!�u�����H
5\A��~~�no]Ն�?{��"���oj�t��Ѭ,(�i�m�X�'�F�!m��a\�/�>��4~���X{!,(�'�����ꤐ���s����%@M�h?����D��D@���P� I�i��^@�4|�y�_=�\�M,�P�&ޗtjM|���2̶ wLQ<��|��g��ORm���	��J}f\[B��U��<R��2�%߹�v��9�������n��k_���t�|�mZ�euє�F�0�QT�.�O|i+ׄD6��P:�p-f��mK)#�~�������2��͙�p2p��{7���C}�/pN��Xc��⦐t����E�h�b�
���H����I�$���F���8j�U��tD���~��m��95]�0v��	��x�D�{�������W&T�1�QI50��gS�-��灀 ��S}v��k� H0�pG���ȟZ�M���>hWt�L�'��T)E�W���0 §�&��C\���Әn b��	�~B�Ah nD�{� x�/&Q�4+H׈�X�����5om�����" r�5L�㹪
�Q�_��{>�Ȱ�d:kb� Eh�l����1��uiΪ�����_jh�E<[V5�����XiO��л�7<g&����8=���pv[��w�I��Y+U���1v�T�죎'����8ޥ(�+RC����a����2����$�����r}+F��'9=�b�}�+o�c0Za��&A�&#1��H��0b���Fc%K"E�☖s�EW:A���K$���9n����`����5�-������k���7~m�m��?*� J� tATi�|�)6�I[��$�Ca��v_;��_z��y���횶.�U��\�5��?m�'B�.i�J��G�Ra4�r��g?20�U����w$����5�;b���P��������e�(\� ��7H+�υ^�q��K�3+a�'�%���9�žЪ��O��nG����ۨ�_��tOa�ti����4e�����W5��k�~̋�U�?��=C>v��`�i�K]���'.�)7�0g����0�A8�0�."���~B=��lwf/�3�0
s��!~Qd|Vu~��h]�
(Ǚv�`I��g�VO��W�6�r��e��mz������{!�4^pY�3��ٳ͍Q��c����/���zZǐ���:���V|�`�Z���Q�~��qu�ȇ�ɷ^T��b �s�i�9X~4sݔC�I�a����%�4�b��O
ޝ��8<���(/�a�o7���fw��L�+o��l:U�	Kz:�I�J��X�N7��wV!�N�-�� �z��3�Ut��*�:���D@����{F�ʎ�p�Š�r8u$^%݃&� ����^����[�%��fר�ˢ_�mA�4g{I(�sY�JЖ4�EC��h-���"�l��/T�Qݘ,�{vi�j"�B'Ջ��+�� �D���J?�|Z�!�&�(eFt8	}&q�	�+[*�G���o�\r�9Aא�#o��J�#�5m'j̗��@�����7��HXOҭf�7�E�8�$��=En�3w�zK� W�u��f9,��؇I��;���I:aE�Se�t[]0�Gl���DD����AvB4�����!���y�̡-�H��I����p���W1��lAPr1�ʑ��B�5�.y.s��=0I��o/�-Zw��[���Z���>L��[-�pYB�я��B���+J��>2�AO�4�z^�l�`�L��ᒍozd�:��S|'Rc�=4�.�h�c��s&b������Wk�}Q ڥ)�qn�`�M���V�q�k�X�j
#�5;�A �0	�M��wF]��(���j	[l�>?lP�"����$M8�/���@1�1�N ~�Lz�H�^��{Wg.ʬq��(J�)E��QCriXdq���@w�k�;v����K{G Y梒��Ӂ�@�Ԧ ��.?�t5[��pM���Ќ�{�?��|T&����)�s1�e0��2�#�i&M��[�Y'��"�D㭊��F�t�'�ߔ_}jqw��[��	A944��ܹ����s%"�>~��>3~I3f9r^ѯ��PJxE7�G1���I��c�ٸ�u�J��)��x��r�m58�k�jvB�3�;%��Z"P)������U=p&06�BH-�[爄;;��M�1��Y���� �qq�_�9���ْq TQ/:;��btk�	�����^&h� bg���5��5���L�B8�UȠZ1�hx:W����aM͌hx})fJcI�ν��N��a��좈.�:{�X��V���ć��!tX�qpH��h�lW�rأ�4�cq�O+`0�w��Lef@\P}t��ik�N��3X@���E%�Ľ��ɝ��~��,�x��L�&7�}���X�e1��
�����A>���N��H2N��O/'vi���������i�gBP���R���K�q���09�:ˇae���	^O�M������p2操iї�d�4hRo�_7��Ga]����<�O��l�5g�Oݹ\�Q.��4�*���E�� ���1)(��ށ6j����jw#M;��X	c�� 65�įƙe�b8!�͹$�_ p�U�n�X�%`d�����'�����*_�<ۦ�2kvNUY�:��p��fP`�-I�� ��/b�\��gf(�LS��8�}C�De��`,��_��G0gL,��)k�>��)Cd%A�x+w�gF%xL��B\Mө!M�X3�� �K�Я;�,to��B�+nJ�m�R��*�*=v�JǾD�bX���'Wj�Yv����EV�c&�����ʧ;H������O�"N��ޢq~����7s
��j%\p�?:�TU	�ΐ�s�7����C��
��_a6���ϳ(a[Ȭl�XF�H�ܒ״�8]vtʁA�6I6\���->�6v@�����ٷ�����&)H���
*�cb��]_�G4�6Ϥ*�Q��_&8&t-?�"J���6�)�1XT��a���~��I�;Bt)0����4����w��$X(ȕ���G��D��;Nbt�����_^n�����R�� /�Z��ˌXu0������0ĕT�u_'�fS�?����y�t�:��DXv�6.�������m��Y��iSP״)҇*Rz
�F���^��̠l�2nUq	/����N�n}���0���H�nF~Ŏޅ���!b� �c�wOZ�7Z"K�{�F0���������t��ZV@�u�Mյ�F��kU�g��]d��ՑR�y�m��a�Qd�)2�������o���0�l+Ҿ[�r�$���N+�y�XA�X�6�4w�w�.��a��E(�<5�V��d]�;IƛY�#Ⱥ7���9����� Q҅��À�;븣�& �/��w4FZ�3<.椧�0�W�oȐ��h�J��>[�5���$1,��I��|�Bȝ�d�,1�?`�t�$W��,w�l.�&7{ػ:����uZʢ�N�_�I�MKc�E,L�6��8d�qؘ��jo��t��L��`���M[~u�2���GT��HIƐԙ!������쁅�s���&Z��lx��!����Ɣ��bT��dj!ykY�\��u?� �b���S����F�U��q���>����Q�@yxVxS=)��_�"��PՆk�I~Uכ���.�%O-f��f2���}k)2��aB����B��gW�Ч�byj���A-+AHN�zMOWӖ{��K};qZ�
��v��ۈTomy[��7�HQ��N+���"4�L��Ï��풷cU�`)-����1\�l��/GE�Z�K�֐c�.i<�I�)��Uጿ
{l��;%x�0�W�׫od���G騣��
�Fy2G��7$v�6����Wm+�x��U����IY�RB��(�(���씹����d'�^N�,	��� ��4qݛұ��HAW��!;l��c9R��-�ڤ8Z'm�n��-z��"�V����!�1�z��������8��ɔp�a!��9�GQ����M��PcO#,���[�}� ��I�/��,��y��(�h��������� "��]Iڨ_ $S�@���IPa�P�� �����s�,��S��imw��}#���*�	f��ڞ5�nE��[��r��l��k��ͦ��2��h�X�k�q���~��:;��U���A�Π����M�h�N��]�<�%#����W)ew��xU:_ [7A%�����m'8ܣg�n���~�F2� ��D�uS��Z.��:@��[�K��^=��\R��M��%���NU�P�h��V87[F����/�j
���uE5$J{I���L�x	(�� uP����#�鍲'���{�X����nG=�P���!>�񻻕[E�8U��#*��<۩^7��\C�ZDTZ��t�k�� �朐4��{~X
0�RY�_bmQa�.�M�F?�,B2���x�a��C���U�0J�_	��F��|�I=o��ia�W�<xSټ��d2�V�`$�;�Mޅ�_>��V�R�W1u��Q=���1��8ʁ�_b�0�T����휄�J;�,�%���敛0~�2	{r�B���IVr3��A�j�41��D-����~)�:�ċ
��`h����H2v֍����\��m��]ĭ띅�u�Hi��(�@%uɧ���3MA�Y5�>T�`�K�F��9����5 �+���u|�>��L������T��F-�7������K�/���a1�K�fӇ�Bv��,�@��}&��a�7�jXB^�o���/�}�<�S���)��KVx�N�kb�V5_�d�:M4&�Nĕ�Dk�|�kۧjAV����S�W�*�>�R�?�������/' �oa:{��S%��1�
͍�9�7b9[�.�z؎f��,o�������%��m�_���G��8Խ��퉹�w��G�_Iۡ���3
T����W�1B첆�jݺ�����d�m({0��B�ݫ~ $[�4�@���5�m�"b-�N�%�xb]�������_�ߐ�~�V�;��`�o�ї*"��t�f,��f����Z5]S����:(�I���X�_O]�. ���,�uƠ�5os\�f�c�da���!]j�ܠ��k�Z8ԽkX�c�O�(�o7�,_����L�T>���nV����3��>xքΙϥ`rj�S�Il�{ѾE�]l#t M��s��T^�Ā�E�!5��%@~/rj�r���x=�J⧻<�S���*Zu2P���+�} <��p@�p����<$�[�Z�����/��*�ۼS;7��an�뼏5��j~
��`E�M�<�d���	���Dy%l�O���l��:k�hY9��WY��u��]�s�B
8��%��#����6�+ų����i�)t#�EX�c$+�|2�[꒧��^ڗ��d���vѸKz����]u̅�`8���SDL���ɲ��DaC_
���q���g�YCV̏�ײ�����_T������g��6^���yT�b���>MS�C�]Ph����Q&�]dd׵�5�o��ƕF:At�����C�3��fy���I���,�&Vܧqv+�X�/D�r���.�i� �V\����I���ͯ*��Մ�i��Q�	��m����=�t�1��6�#�,��]5���d��f�7H4�߯�h��w�B���;8c��N���N��C��2h�ݦ[ym�+Ǿ0 Z��`����53�4}��������mQ����-n�N�x�դK�"�dS�b�*˓�L���q������+�D�Bv ����V�¶	�`��K5���4�g|)�� S�7NN���Oٖ�7}�}�җ*']���]�����,�^@@yU���)�(��^��}�DS@���%>�}�g����J. ��X�+�R��	EZ�5������Ct���S�GT�H��/N���v�Ml�����q��ŷz�l�<8#��9�LUb�	��$uἂ�`|�	��mPVXQUp:;�8x�d���_�����IZ�o8�oDT���"`�&�������!ff�ʖ�����m�~�T{�:=��S6��D{�r��:�����L�K�vq�ٷ,�>bn���=� ��j�0�L���O�y�ؿ�6��i4b--\j�4r�7�k����g$ya�i<bAAް�����k��OΛQ�B�t�M�[�Y�u�uA:����(��v��OS2�v�-�&.����]�ra�.X|�0O6]ٰ�"Il����y���F��[F��S ���*�FQڌJ]ɪD����e '�	u�Se�J�ĨO$��Ԇz�g$���b�z�}�u��ӥ�׬�V��CB��0x��;,�Qt@ڢx�sN`���6�L������������� �����9����0�?�m�!����愈��/���3jՐ1���gP����q ����S]�'�)SѦ[g��N=I<�!<�#i{۞���Tg80���� �")�m�
f��榫�X%���{��&ڬs��6"�꽁Ե��؀kn�j�5-2<��gA���b"���E	d�zpBQ��R�����2�ؙW*�����׾�k��J����ڢ�~~_����96�
�~�I'!���v�@PՎ*W1�/P�E|ù��:�����B�R�\PC��58�'e�l7��Վ�k�Fj����t�sH�;��nWS5iM�+��7E彜4)�` ���X��v�� '�1��������.L��S<��UK����B���+�=���D��~�2�]+���r~�y��f��o��������.���⡔�Dy��y�E�����W*����5�5���_�Z���a|�?8@�~T�~����qu	�����c����
���σ���o�33竜�12����)<�@4L(�����2��	.x���B�J��G틒�dni���h��$uU���IIKޮ0M����X�-���g�@���-]�i�C�s�	�L�0��B³~��Ĩ����BK3��bE��$���a����[�4Ά�(�97�k�i
�w	���?X3���^�J?�J�a�c���6�2-k���,���4�����PyC���e�r&�l��p��B��Buƍ�
�ejtܞ�ФV�d'�F�z�z�錴D�5�#�)��z�I��4rp˰��/r�E�b��P���'���z,
֦��|}�o�8$NϿ���N��X^u���#�4ߌ�j�j`��g�bl]d�	.�)B:͢�r?����?c��|!�q� p���@��\�d����,h搭��tr#hc ��^n��kb�'���i��7��ҿ�q����!�	Bp%0n�� ����"�o�L�����}���q2uM��<���:'�m6a�E���IgAt�6���5�
������cK�����5֜?�"�N��M9�ha>�B�}���y~���J}p���.�wS�I��߶�� LUZ��|&���Ƶh~K���;G ��C�N�S��L���r�o�"8�A��}`t���6[�|$6�S	��!�S�� �S.�}�[k�;��8�BSU+p(��:2:�}�B�2@�Q��k[>�(釛�{��@*+o8�/��ʔ#�y��^�.^y-b��Gkx�b���0Yp�8�6�i<o�P���a���۩#m�o���X3�����3�=E�38�H�"\"2F�d̻sX���[ L�rՂi��ǈ���|��S����S6��1s1����|��f�%���^��:V���O��u�bxЃ���0X���\˪ oN_�O(�X�DA8w���I�ɯa��boxP����1rW���t���ae��?�<��s	�2̄Q�/��SN���o�0��r#c�Ԉ�"9s���]��
Y&t�ڋ�3�,���X��\�o�'_�K�=�`j�^'*�X��J��[�����"���Qpm���$�/=�Lop��b�2�Z���:W��7�	�eR��3}OSZ�a��CBw0�v'���d#��U3QP%q�n�6H]r�.�pM���0��f AON)��,M�	��\)�?a�Hc�aH��٢�'^e�L���-	j�`:�C�Q�����o��_��_���a�Į{E��cP�pF,�.�����n��_�G�mUg��s�w���W9�)��o~�����ʳ}���*M�gG-X���ӷ�A^�}�E��g�B����W�\��4�i	��9����=	Z[��?;�����	�y�0������6 �}�_P��b4�0Hf,6�S��$�55C�&��4V͠ �2D��\�N���Y�c-�|�I`%� Z��/GY����p�'�MNv`�n�--Ur���+4��%�ڎ�^��#�b�U���I���j�Eh��m�2"��i(�#��R
���� '[����"*� �FWZ`�S4W(���@&�X�*�]�C$������}Uյs���
Ԋ0N�+F\ǈ�����?Aҫ�t�?%rK�R��c�)���O��MX��>M��85hҪ�y�VƁD�C?1)=F$��t��I3H�(yE���0��)�r������v���� �T�����=+�\�x�	L�
~�(���4�,V�O'�Ζ�I�gΨ��PZ�OI�;����=��z1�W������!��H�vFP�j�* �m����Vtn�L���&�G!SC�H�Կ+$2]��s�N1�.]ݟ��t"/Ƨխ!Q	�g>\�4b@<��p%��A�����_��άC��T�3�?�֒8��� ���7@�Al����<�c���D�YŒ_ 21M�o��q�G�>�=ӕ�'|�,,4��Q�e�R�,tF���x8b���stcoQ�F`-w����`a����g"q#��~��n�"�
��V�z(�`�:F���(H��^\��A�<�doq�y'!�q)��B^H���>O�ݱ,�cd�tc�'����#)U�ˮ�@,K��a�5����w~��������]��?�eZR7���y��S��\v/\;�EFxE	,�Gw]�:�c�+�Q�(�
3�ަd��lkY��4c �����?��&{��	�Oe�x��d��82b��£k��
�
��ԾE�M��O$jAl���W��'�DGN�x������u��m~�2e�0�t`��(xD������h"�+?��Qɬ�ȹ���y��y��Y竇���i@��V^Nx���n�3�z�˦�|��B+��k��h�ƒH�Z^OM���ZgQ߭Ӕ5c2��5K��g�)N��K���M�㒱�u���j�8᫟��8�M6[}ƤT��s�[��B��*��T�Dmm���_�?���6�E��)�|��gw��ԥ�W��`z��3��Ӿ�8�2ĉ�G���gD���ЁO��[���иU���y��.F�����)[%�x���0�2R�$@�Dg�\S.'p+��_�H���|_1ؘs�cV�2H��
����P��]K𢐫D��q��ࡅf�I&�8�>Վ��5���T�~����_碩��T�#KrR�'�Y�3_��¥�N�W�Y��E��]���H�9��ƴ!���ۢ�4�-�)�/�W7����-��NA�pZ=���v�H#h�*��|Haj7�N�?��B�.�`��F�҄_cZ���	yH2�`���Ó��k �����tNx*EZ\��iE�w�7�a�^�@�*�(���n��'�htV!>�!;��z!�ő>�9�л�6(:T��}�P����	��(3h�����L����
������j��W�����#�]W"�ݦJ�@cYf���i��v���\;�Hc���N�&&-��a*<K�+�m���
<�" y�Q�h,�����	����A����r:ř�o�8"]R��^i�O�D���7k�����ּG�ܲ|Xn��w��2�}h�昭㳈��{�V8�s�-�
T��M}Dź�3���� ?ԍq�B��NX1�+�m���S�����'���TD�mx����!k�q=!*o�f)����J�gP�ʛ<��������(g��øǗ�I�I5�%³�NL���>"�gx�����r�c !�'-s�_$���8lNO���> �7Y�9�����)$�CW�r�.���W�s�t�H�ܠ����
�S���=��C3�mR����S����|z~G.�#�Tc�^����+
uC	�UO��n���z�G��#Ru#�R|�3/c�KӐrP����t`�S�m6zS�D��sK�mjb��>a��,�K������a��"C]�p�Tgi��N½Y�%uvغ(F7��Y��bN�D�7Z�!�V4#~	�.Ʋ 
�O��>�u��%g<xO��7ȋn	�궙:�l�Ǥs�#�����l�Uc��w$K1�4��Z�F��L��{��&��g�)!c���V�O�I}��z�An�z��I��|�s�!hN��_!���0^�!�嵈�~x�I����ZS�F�6���/q�`#J��:@Pa�+TR��Xv2F��D� �2ݰ��������Q�V��0�_G���C<�k2dn�0��\d*Ȝ��^R���1G���5>r��	 E$�D��V�q��V��B�������#�D�C��/��B��Omq];����c�z�Uۧ�ȸs��e=�̾9�<���'٤'�\䲎jw�5FR!�SU�3fc��г*�̲@��YH�����_�Sm:A�xX2�զ:�9�-A)>n^h��|}���K%'\���mMW/
��{28�=B�/Sc���R�����xc\5����bTb�l_j��[c�J�%Ti%O.T��&����b=��.��A���}1�ʻ=$��"���n��*��Ȥ���((8ƍ.�$�xT$��1<����޾������4����=t�RZ�8O�M�u�d?螸c�Ⱦ��ŵln}?	>��.p�PL������`��M�[ �B\��٥f�U��I�t�^hg�Bu�&'��@�^*��7#��H��Ō�k��Z^�B>fDg��)��DtC͈�X��c)^�nc���/�9WyJ�t�f,��z�ⵕ�8�j�����q4MZ!��ȻR}�xq�Db��d�fѽ�_v�[o�ӶZ��o�,J���7ȕ<��GNd!�قI��{]|oD����H���7(�b�{nAy��W`�HD�9���2( /��4��1ū"P��XN�<<��@� '�IU,;�P�N��=9\3�+E�����O��ܩ�H��2ԂŬs�@�i��l���n���=��C��׿��4X���bph]'���o9�r�Y^_�̋�IE�M������.'���r��&�"�e���cK���}�GMZ��?P��]����3m.ӽ7���B��{T�;d�X�~���F|&�C*���T����fEۙ����1W���0�wvؐ)f�=^� ��c�`@G�9KF1�[�-�m���RA�7=t�?�ψ�yB�^5+C����[4�����X�s��-qΠ�#����㙭?�w��Q�؉K2�O���R;K�c��+E�{���=A�����RyK�������@��Ui�vX`�Z����HI����a~�S��r�~��y|�r�"?1��Kԅ�A�8,(�fr��`
*�X�Z��Y.}<?����R���hnc=�5J�����k-��rFg���/�e��1f�H�bAF����d���lxn+g��n�ح�y�J�լ�4����A����Y�1t98;��_����dF|�fF���8���ʷSCtG%���XY���v�C
�K�J#[�ϤR��Bֱ�b�ș}c���t$<���S�d1 2�/�ꞳY�_�2�4����	8N��X��</c-�����r �?�06|I��r�u7��­B&{�	�Uu��6��ٔ��� Q�81v�c�׃��tm�v�3�x���ߗ!IK�����K0�~�yc+��^�kKf��
n��4�3y����)��\)b���V�Oq݄��XR�B�Q�ǫ��G������8I�\�<1  e���XV��3~�����NWo��0��+�k\$�K�U����Q:|CK���V�r�ǹ��2M+�~G_���X 	U}��]ۃ<c��p�+��s�7�)��q��Z��NV=��8+�y�n=�xzr�W�s�T��?dݯ�B���К�k��ۻ�36�J��((����8����Y�S�#g���54.�.�����Gm� wm����en��8 R��Jҥ�o�B���y>:�7�i(�' Z��~DZ����"�KRB���� 8��[�BU]?ʐ4K�@�Vi��).�,�������|�Xs+Ń��{�[��٫p7�:hژ9lܫ�(9����i=���v �u�l���
�}�=��z6�k�&������0,۝n`�f�4]\ׅ�O���vA�~��l�q�D�R��k�#�2��%Z��	������\7p��J�|mu���Ӈu�/�O��5���,�^���N]{)�c���O�Kx4�#A���?)���6 ����儂pY�S�?��ڍ�>�8��i�Fսz���`��a3���3���o�OV����Ǩ�,q��Ă꽖�)��I�$7����Q/]W٤z�>�8e��Y6�Y�T��T�'V2B5��Z;r���0��'�@��*;Q�����y:kW�����RL�ս�wAY��Ŧb�-|��&y���<Puyp�~]���g�;��J��x���ti��kV�/}~#��BVIɮ�c������3ch(y�z8+km7b8�(0��sb����0�d^���%�߷�s#/����=�KX��(y�y��Z��}E�;���׹	�x���Ҧ�e{,:6M71S)b�~3.�Ew��<�%]�j��:�:�z���E�����&�F�Sӥ!���0U>OK��V���ɪ�u�-�����ZMo�"�aI�G'�.�E�=���1�I��*dA�y��5��7]52"#3t�h��k����A���$L�?su��W6{hc����19e/�hS�t���I�k�����d�KZ�Q�vl���ʾ�;L��oN�6�W*t��� ��)�w����U~�dM�w����T%j��Eٓ_�KE�@$�咶�v/q̼��e��m)��:�c3ay��L���Q��M�>�����N;A����q�N����EVW⿬�s��/�􈡵�\����#��o)���b|~�jR���
�4�lb3��ft|���(���!��_�&@Oz��Ge=jU&�*�X=�U��kC8�U޸!� ���8:��?4э��S�SK �ѩd?]z��w_�Rh�����l/�{�	�-
ՙ�p�Ͻ�3O�+^������!hS �=<C@�M׾���/�j��%���M,��+��D��4�W���s�z0=%���P���J�
\V+� �5exz�E�o�ڬG~ѳ�j�m�,S=�d?!C�7�y�ν|�w�	k����I ���PJ�D��4>LV*1������^��6�1C��b�3�Ü_r�&Q�\]�Rq�tT$u�گ݉�UF^}U�����6#C6޼������`߶�K����R-�q��F4=HO����[{p���z/�=P��%g"�H�!!��8�M���Ư&�9��5�[_��	i.�Iڲ��#������U3*k�����	���\m�R$��Oz�W�搀������^mg��ˮ<퇏^�<e��懍?�z�tXJ��,�C_���c��`#���[����x6�n���M@�7�V���[֖�r����'L��>����.K򻛗w�n8L�.�H����w�>|ʦ~ϊ��xP�cz����!�3��*b���]�N��#S�{{�\+�i��Q&��\���zpF`ݎ���?��W��4ì�ךN��i\��V�����}��ډ)栜K�����2{-�)��BaV��_!Yy[4Њ�Q��7�p�V���Ω�;�N��:��ec̵�k��Xc^(!���ʹ�`2,M"ʥ�v7�E�쀙���JSnM[���6�M,�w�q�����Itoq�Ӓ���5�M�Vu�U�����8x�9���$� ��E�UI�]5`���ش��.L�o� $��5b���2="���_����ff���2Un[ ����$w5*�r�>�*�x}j� g>6�]�[z(�;�E�+�~����t�H���}Z����4��?�P���H�l�K��}�J��>xn��G�6)
�a�	����'5�O	Y���X/�������)�x���r=c�PG�]!j8�I��X�cƒ���K�R������cW���lk���sI�މ��Foۦ�E^5��4t�/��r"ȊB&�Q:��x���sA<�z!�5�OYYHa tw�G?��v缍-TGS�1T/��F�������� �O��H���n��is��S��zV�I��ͤ����q�=G��SQ�T\���8��ϱ2�?f0/Z����N��18b��+"$C��ֺ�p��l���Uǫ�8
!n����Z���3��6(�J*���#C�:vrܗ�H�}��m���Ť2��lX��O����`OD����""SI��ȼ�w�"���K��+5{_�����d5b��,m٧���[��7��F,�'����-�h�+~&��5ɌCК'����e�l�cv��s�{�ifrYiK'E�ӈ���E>%f&�ʘ��TP��,6b揅��lץ�����oa<�����V�_����gW���$��W���E*���kn�#��-���+��j��g���4�G3�#D�w�j:�w��uU������� �i�v��� � T,�+�+Ej"<x��ٷ�p���2
�D��dG�9~�R���Ʒ�<>t#�?�$��y#�j�}H���s]zsO���]�߆�.��x��]R����'�0�e��!ݗ��3k�0nӎ���&�lZ���ݼPa���#P��jŰ�@�z�"�*`��-��'�P�v&Y3�sq��BZ��*��z)��û"��:����`��V��H�RC��	Zv�N������BA���Ֆ{�3HI�z�������L�l��'j�ٰѱ���!�9�6�=�B�bnW�J3�����yQ���]˓����e��|;�gGg�Ĳ~
m�1+�UZ�Uuމ9���nM����rl���g�yaӸ@|�h	2����\�JdtG�3��X_ؿl3��;�w���@��\������K5t<�"ʈ3s.Z��7E�W��X�m��쁗Ͼ��pg3���-1H����-���ؙZ2��?���t�X���A���&a�l�Y�z�Ϥ�B[�}J�~f��LG�;:�C_�<�Y�����_�*��r�E]g��Uy��G,�R �����~ɶ+ ������rk,s�M�%ib�^�wwH}�v�[� �OD�|�l�p""��5$rtJ�=��k�K�'ߘ_'��j�I��6#K?ڨ*��l��O�N���m\�B����h)������9��
Br��
K�iA�c�$#������h�-q����<�fb	
�]?W�w�ƚ�	Et��}ߩ|�:V�[:O��xM9��l�l�o%�]�*֕��܈a�����~�����jFv��+ϴJ�{�~���ݻY�+7�J�I"!dn>�V�-�P�T�	�93M�N�'vAD{��&Vm�V��=�K��"����NƊ��W�[L���K���%g�7��h"�Bؾ��F^�j:��y��l�f#ϲY��A�ơ��j'�_2<�H�KxYPT�j!�rYӓ�*�����l�j	����WQ�S���yP�~-Z�7d��K:g̱ʶ-�7`U&�d��%��o������jM�I@өH���1T��{��rF*�'�ŕ�G��.�?WK�ߋ��:�ey�{��p@�F�E�mg��D�#@V_��R1�^T�����y���x���-$���]�:��C�ܟp��h�yp�v_RKb��O��܉���i�a� �S�����c�@�摵�
��l�%3d!33�j��H�q6P�o�d�Еb���:��c�8���@�쫹��diR����<��B�J��ZX�}l�bX%�BZ�&
ˮ���/�R=�u>R'!��bE1��);HP�BS���@Z��=���;����4B~l?��� ��@��5,�W��2�Cx�!��7�H,2�nb�	�Z���oĦ)Վe=�@{ K5�@.HF�0�`��O��(���)Ì��K۠x�H+�Vx�����=��nL��4{m�ǭu�"�&�^=cb@?H�����RI
�6�d�����g�M�w.�k��ΌGqb�]�lF	=e�k�7ryQ(�'�7����J9��wt6	�q�s���p	$��������g��i"�JRN��Qd���6cї�w�TXr΁؋�Nt;5]?qF OH&�ԕ�ww�k1N����9�΁�r�������Z� �����s�J܅\{lo`#,�ڀcBHG�n�ӓ��A������O
������yw�w	;i�����#����n��"�!@>��k�x�4iN�\��Ae�܎����˹����	���TE荟1��T0�U�:;_��T����oH#�Z���8I�d#��� ¿�*P�JD-Ȃ���S6�*�A�w��q�1���r��)��������:�Z�(֔z,N�r�Nr�ArZ�[i3;i�Ix�lWs�<����}��98E��:zM�W����Z	�"�-*�j�g�J���߳�W����h��S�Q��)�g�]q��Pv�05������׊�87�ꈹ�($�I���Z�գ�����'m]i�J '��Ǘ@ɽ�����-��?@�"Z|�ǧ�m�Tڸ.X�9K`��^�v����� T��<KS�*�ujΏR�$;����;��d�`
u�6�3x6b�h����y��ı�|��P¶�\oD�wǋ���zÇ��Q��e�h!���	�$ �G�໪Eݎ�����z��]w5Yl��5m��JlL��J�<��M���og���c����L����̢����~�
k5�4@�|Ĩ���5�	��e*�88(�6��q���0��#�?���U��?����\܀��&�b���,[��#�Y87�#e�|A� DR��N"�{������;�B�^�rKu84�~9X@�J@�q�y��P�?�z9MJ&<��]=�L�.��ױ/>&�� LnD�i�2��Ov
B.�j�XM�(�"���r)��DI4'��Y���|��T���B�Q��W�Wۮjh�D�(��H�z�#!�;��`WBq�g��؇-�{aP��P¾����Kj�ے��
nc���[�c�k)Ս$ؿ�\<@�#Q���x�4Ω兎�NU�����)����
B�`�oBe��CހB�&>5�W)"$�r
�?�C��D{��x!,hT����D<�R�&$��q�u�7���YanU�G�[��	��3��8�[s$c��Ń�����n�����.�e;�C%W�7��;qs�Ҵ"��g��="�ѱ'1�ۨY�
��]�^g�V%*���P^�Q�7�L�Wf���a�z[�z�RD����<�be�$�Q׼C�Ґ�x+bwڐ@1�87���b��S�k�4��k��gՖ�,���t��R�ֽS>�G��+�4���%��i�b8�k'#�Ņ����q_pv;L`)-�qE�s��P�(4m�ǻ�[F�D��pq�q;��.��\᰻��b���7q��Eh,�Rϭ��c:���f��\Dٯ��U�i�����8�m��]~��c�l\i�	�-mZ(����/@τM}ð��S�u���Ұ�1�M�	���k�CZ��e�k䥔�����
�V����kR�Y{�w�W]f�xq,Rڭy����6tD:.u����Cqy�=`�����5�i�,���n� BG3.z(��|fj#q�z�f�8.2�&�����(�;�~���T��S�1�_����	�JQ�p;l���Nk�2��1��W��awz�a����3ܚP	��/�Fq�l�ƍBHQr�ў��M�A?���C� .T���V�?�6�Yń�S�Daq�N�?������n�`�CQ��z^	o��t&1��:,�x�SA��s_�)�vt�&�	�Rt�-�4��/!���V9h�H���'�d��x-��ͩ^����xH�C+��*x����N�}���'�͡�P�
��&���c� ����n�_d����5�#�Wt�L��{�//&��P�$��|��ѣ�X���.��B ���	�u�N0��V7z|��]،g%(���G�p*�}�L�@�%B��t�;�����a0+�e�`�;���飃Qh�)㘢�����3��2T��q@Ѹ��2�fz*'���oEIh"��j�	�|4o��5��K�\Y�L�$�]�&�Ti�j@=��}�=;ʞ�/�0UN��p��k9��K"iK����ְ<�C �Q;�6q<9�KW���牮¤�`<hX��@�8��mȲqL�Z���r�!������,x��4�x�\��N�� jc�݋�8��kD�WM��R�ᄑ,kX7�)b���D�OY���O��}��vLzW�K]��m�Br�h�Luiۆ�Ws=��R��&��х<dN0�5	�9�z�_W؃��!B~�	�~�d��(TaQkx�4�� yo�/KM�K��'̛�S-����b�YHZ���=�8�,�"h����J��������(�ClD�$��I�#;�*wO��-D��1׿}+��9�@�\Z�n�r6�>��#�T�YW@��o����o�1���5�j�����ÃK�{�mQ� �L����T5�M�I?6���m��,��n�6�����BU��B�h����Z��	>%����̳g�B?JǸ|7[@rW��!���Ѵ�@~����'(`/XӠo�.��U^7�2��(�D��-V����P7�	��G@z�/��*X�W�<�w��c����Y'p��I��K���\Ln��e��r,�4����#������oDǐ4�aC����Js�{4���%/���>D����Ų@�4M����%W���}h�T	1
mΧ
�x�>� ���;l�4��R���S<��ƹ�bTW�նOD����L:;���H�c 
�\�������[wC��Vb���a��v�z����ǫ+�n�޻�$�pR�bSb�32�Y��m4z	�/�Y�F�p�G��������(��,N�{S�M�#�u�CGic4��RG�u�E6�5��j+�,�~��\��9�j4�e�c��﹨��-��f/%;�����'���VX����F�e;i.�<�H��_-8̦Z�K?H*k)5eCB춛<و7��K�l���-�(LW�L"�]O���[!�*�z���C�T�Uy�x�s�J��P:�r��p&�F��*܄���)��x�R����x��U�d6h��خh�'3���/�T���"(�d��Ohߪ{UE����KBs��Z25S�ܤ�� !���-~��o){��G	�Xňuk�<�C�T�^�T��n�e�tN{��ٻ�8�yDz��M�I v���7�F�O��4s���ϝ~z���ܮT��{�;����y�eH/�XMAg;*��2�\�.�����sD��]�T�Lw��Z+ּ۱�ߠ��x����� 3�/̾`�O�i�C.����ݢ5Y\o�Y�='"R5�*ğ"�%t�wڻo������f�a�99�X��׺z!��̈́�I�����޸�<�S�ZZхVb[��ċ��`�Y���Z��;�s�._�j͂�n)b�Ҿ����J�:���T��޻j�����w?��eu�Đ�cHx�3��6���̾un m��u��q�L�	�ڲ��M����d<��Ռ,��������*�jSU���c���!�P2��}�Z!�A����~=���=$�S�k<�v��T\j��i�lb����K��fL�06\��e�� �a�&�11�����r��# ���|?�"3k�G�Y�AM��8����v��9/ 	���W������ޢ���7<��6u�ɦ2�L��򛾁c���5���=FQr�5:���=!���ô ~O�-����Gi[|fm�|N��g��WME��"�����(=n
c���	�e�C]ǾV�1ͱ���[� ��`�z��V�ּ@H�a�ߴS�'6nq9 ��L�dƻ!'[沙 �zw=���f@:[�gn�YyN5G`����,�����nDm��ej&L���W��q(�4M�q3���LA`��)ufɄ%�6��%7 瘛�sJ����v�!�Y�s�? �kV�(=��FSM3_��w>5^VW!"9�	T*��\��|"���iF�:��0>�_v"���^G.�c�YV��#��3��4W���)+oQ�
�6+����9�č
r���$�S���"��r-�ёޠ�=�D��F7hy^O82AF��1�����l|F ��3Pl��o+���LiX`
Ds�꜃Jw��aF#k�x���)W1��\�$����p4����Ze��_��R�MA�ET���@+"����.����J�`�D����3� *�PՉ��0�<��$�߅.���AI�b���h���
ǃ�Y@p0Su"�bf��(�,�Z?|��F܊;!�%��Qx;� g8G�7R�'U�db�+T3�q���m�!�	�! ցۀ`غ��饸/��n��3��$���r���f��Zm�zsj���Z˹�JP��y
oR2���a�*ԇ�dg5,MsZ�"���,P�{)�y��Ru����i�m���r~�U��n}�Μ�z�R=)���0#���{	6�G
���C{	�"Nv�Ʌ�,ص >�ͺ��2�*/��l����WK�@[Q.&֧1�6�����)f�(~��������3ܸ|���z�[�l%i#�+�`Ջ���)n�Tw�xƔ�"�ƒ#:�c8�5F�@fz�,�z�"@sm�ߨ/�j&�$r�#�Q'�m��=�v��oK,���?�r�����qK�z�C�٧#�pmT{t���/�q��)��uf� \��~�p8�U\X([���%x��L6�*�����n�b�G��������&-��m�@�j.cT��" ,����m�.9�T7Sųn�ap��=� �"�.懳�rLh��uj�m�k�<��f2k�ħ_p�(w��� ��b$O)�F�S � .�ȡB�eh�%�1�C/��C�f@��^;�Z�Xmy�.�&f�"�ɥ_L�ɗg�l�鸿Ny�^C��>��^_XFjoM�e[u^N�@���'+C��+F�gQ� ��Kjp�0��Q���1I`^n?s������(\�s��9X�+Byb8a���P6�7��~��"ͯ�ױ�.����Ղ��Q��+�5�������?mJ[q�jW�%Ԩ$��$PV��&1K=OЅ�lm������Ϯ��$/^P�h~�#I���:,I.D�R���:+����j�M�����O2� 䅻J��������`Y�1���8����Y�w8T+��.����&/E&��U��E��>I�^9MZ���e]��Rw�ӝ���U��X1�є�����L�b{��r���~+��&�%��sQ�4�-�\H�T����0K!Z<P����;�pz�]�L_���ي�O�R!=n5�;z�o��ڐ8��� N�/#���;����`��/���T���Y�
jL���ku*>���-�!G��v�0RC���4��@9U|��=�?�}����b�!B�*|lw�V�׼�m,c����'�����<V��]o4�SnBv�R�Ib5�>(���,�X�6V��޸��ð��3���У{9Q@g����4H�@2��a�(��XE���U�^P���W ������d�O��M�J;��*�Cn�>g�.h�M��jw�L��yn���T,�N�Ҏ�a� �L����.s#���D6cث:��ظ�c*t��[��/�uL1��K�u�`��Cc��"9!~.��](駰j��=(g��E�����+Pd����j��4�6�Q��g��^�/�բA2[�����)ä��M�r��M�����j�/���'ΝL5i(�*Yk��X�,޾8/g�)J�C6���ͻ����h¹1�?d�o��fa'ѩzճa)���Ш��Y; g#)��gT��Q߅j�29+F N�Fˤ�ii.�1�u��J�d�JP�n{�Bu
2�f�Ɠc��`9��9����6�h�y���H7�g��*4�@7�t�-��b>�@ ǥM��F#�ϳb�vc,���?���1�BxeZ��_&7���U��	��:�3�S3��Rr��&���m�bd����L{������w��I�:�5���
�,�ލ�궀�t�� 8�hr�?M�� FZ�)$4�FX��*�p��Y�4���M��E�d02ؔ��F�d�31� �b��U0�;�_˒џ<QP-Mvٴ;�p�=�?���4&wVj��Ts��Rb@�"�����.����+�[	��u&��f���v<���/��'�/k��i���7~��]��,�m�'�:�5RϷ���?��L��n�#�3���T0w�q6��_����06�҇^��L﷬��c��}��Wa�B���#�ۙOd"��<׈������8W��
�,���Kb��YF�;�N�ir��4�yQ�}3J�Hӆr�Ť*���g��ZfE2����8�]�޼�3)a�ž��i�2-��������z���YMت�$�P/_���B��VaPpR'񜠢Q1�C Msy��O��;L�F���J���^�^ʲ�)���-�������~+e-7�ف��Ua�_�:!$�"��(����,c�cщ,���p�=Ȇ��WqT���;� M֞zA�("�V�F�Q&��H�jʼ��Au �J!ѯ����:���TA,�
R�C�@qs_��7���Ւ
���!��Sd���z�B�>f����֩X�Eo��rK��LU�d4&9+1�d�K��J��Hc�Wy�3Q�>��_��O�`j�cC-&O��a�yVx�l|˟��_�b��`cLl�d.-��&�Q�v�}ݮ�м�������=�?bM���z5�a�7��.o����<B·�|��7����n�u�`*��
�p�IP�p�)c���B;Ç�O��<� �}��L%uDv;?h�"{`��Oag	�'�4�"Ǌ_4�c�l�5	V0M5����s�_��p@�"�`���r�������V��f	���C���o��������O�]��kD�w�C56@4�J��E�͙�޺:��{�����ϮL�4a��ZP�r�uE_�7� !��> �\�!g&pT��Hu��.l�xB �_и�Ku��Q���%�tuVKtސ#��(�a�$��&[�X����)��
1�<�h����ƿ�*t'ժ�Bl�#�b�Cb����Ҙ�y|L9���Y?�c��E)<�����9J_HWF�^���}�)�dkş緔!�1�vTē_�US���iW�T�h�?,����)�­:#��aB�����X��J9��[ke�=Z�#&���B�X��XX�_q��"Y L����V������"�>�?��\����՚�̾�G-�E��{�^��m��x�Sc��7hG$��>��D�(?~�{j��`>���o�khDG}g���pTzJ+3E�6�Ϻ��V�@�ۖ�}[9��1�0,*XV#�O-�>�l�K�9-��k4��d/���+7^�_�7`\�����&t��Tf�U�(���
?��z� Ǧ3.���J�'��!7�=��a��
�2JM���n3�@����g뚯"�$��F��<�����D� ����I���K}�`�{"V��i�#��C]�jh���Bl5�~����h=c��ش=� ���=0��J��-�0?�S�3�2Eĥ����D���$W雗�@��b����7r��x�D���E�\t�����"�ٝ��y���5�O��R�?ě�ʲ�흲���j������+��&7����+e�q����u�H���M��W K�ؐ)m�(�4�&�ȥ,g�:��Ѣ��t�Ha��5�{�~�Y&*�TT�܌ �l��Aʿ�$A�MeQa-d�>��:��l��B�s9���̆C]���Q�q�ŢX}Ÿ�צB�O�3,OR̙}e��NVɜi�����kR�3��RʘC�(�gX'���f䟑&G����<�{�E�a�Tu�>��,�T��*���EF%��^(0��Ŕ,�1Cz�rs�_!4,*1(B��](p��3���G9ĞRNaH|,B�.��*��Tk��}
q�'�bC��Rc�J�Y;�oΆ(ʤ����B�:��5��j�Л]&�v`�p7\�w$_�y�`C�q�\F��\QVU�Q�'�|b���V��>*�A?1S髒��s*�� Era�4��[�4��	��oO�v���mJ�{~:�O
q�C��.$N���\�gD�\U��6{hZ+��M*���?����S"̤Z��V�k@��q&8���7X� *�ް���Z] :����@=Oq�"~�l����
U��0���N�*Ǖ/'F��+X ť�LZ��ww��]�����طEW�\
4�a�*̃i=�8�S��I� s-�������nTf��|��(�n32E.Z�ץ�D�6�N��nXjA���݁B�~p�0��L`I�>�B!$��M�(]K��X0��յ,�b�"g��ټ��D��4��R�H����^����X
��;"SG�&z��P^���]�R>���|�ZqƤ^5�Ba��+�ӯ���)d����b��Ss��Q�B����y�Y�dܡTS���-�߲�k�)Nm��b~����W[�0ae��F���S��)�[�o5�#<��⋿+�q��_�G�逳�@qhp��Sl��UW��i�e�,��igj�H�Mr.�:�`۾;�'�35��?�h!_�ڬ�U�S��)D��ٱ-���;Tҍ�ˉ;���=G�w!_�aI�~�r�ũ-j&à&�1�ǲT�û���T�ץ�!�N y�e���a>��ʖY����g��x�E��.+�2�n� @ڔ��Pm��Sq��S�hZr����e���;^k�gKPC
��=�=�VEw�uk��ѣ!Y�f�����!����b�C,��Hn�[M`-]�@��̥9c>�9f��X�RV�Butwj�,�0�n"l޸9��w��z�'�g��r����FE�}��[��@�.q�M�F���q@�O²�x�;o�Y����:�2�j �]�ڶ���s�BW�����s��󺉡)��^D�-h�����i#�9��Aw��˃R�-Z��j�����Y�|ۏ(�Z7M�d0�q]���Ӱe����(0O�=�D���?U��YwUmV�>��㗀�wh�3��2�i{���/}�ސ�C����=�;��ՖTR=����].s� ��r�HC.�	16K(�:�c���m��.ޒy�O�RMо=��J}�J�Ϫ�6��������)���Q�r�q,��nɅ��;`)Pnt�"�~-�׏��5k���I�J�8��qW�d'�����s9�P�����Z�u6%$x|��P�zx�`ێ)�9D:l�}S9e���V"�jv��b�_c�2�k:�|�'C���k�Jr�"^��'9�c�m�P�"U��"LM�v$��7v�#LΎ4^�D?�1�l�/ټ"u��0q_u��F�'�����E�l�c�d`=�%q�d���p3��[i;}	;O����b�4NQSR)��	��rt�6 DkV��i�
�z�'vKH
>�xlUl��ɜY��),Ôb���@�����{*��j0ŧ����0(]��Ĳ�>�9�7Tg�-�WҝT{���]���W蹱L���D�Ǟ�A�"Ҡf�lY��q2xYm�A�I�|!`�B+Kt��Y�醘�B�ۺ��_��?6C�B{��P���aA��r��[�>�=3�8�ӋsAx0�Mjq�t�jֶ`V��30G&�B����
/��(�q��5[}b����`ߍ��H{��{��n0&�R��{����0�n���_�0�Λ��[�7/��0U#�jXwi��J'���.�lY���5a�/��f$9G\d˱�Mp��v�P�>j)�(XI�����E0���G�Zq��W�uM����rt���A�����NY��r\���/�j��9w�Z�j�"v��j�W-]Y���]������-���`K�!=�J(��;G�0���&�7E���.��h����BA�`�/?��,~��x*mV��5 x�-�,u%8p�)�GE8���~�}����'�&;�"qa���O�8��5G[u���t��p�3"��IƑ����ZC�^�ڤB~�SȧM* �Ka�PI��h@-3����^A�Q8T����k�b�	<����O��,�%�D�`KD��^��d\�;��P"|t��@~o��싗��b[�փ^Mu#��1��
A6#����o'�9�4Mn�p�����ɦ�ιN��h1��s2=��&��0C� ��*%]������ik'��0U�YXjo�G������ &T��Ωz��L�q���/�Ap9;D=�����OO^�M*.Te��f��_��,�{�B�YE&[G6Yo�����L�^�s�����eE�xs~��եN<4�)�{MQ�'�\V��7�ɶZ�ǸP��F:$W}�/��Yy>"���!��!F�#����D���]�]�Y<Ći]�9ٟg<�3�z���+Me��^��K�= ~����T~������"�n��]���WK�B�ҭ��g1]W��G���2MS�å=4���F����A�����j�E<�� =`3�Ԁ{����:N�]������X�\�Ӭ��U$�F�{�DgOENHz���=O��Ⱦ%X%�) 
�V䚱�9�v��J�dC&EcB.�if�����<����6"2��y��\�I��� #����h]un� �oQe?��7���;�SHL����I�0�R�߯g��W����>	ʪg��ueN�*����.#i��ѧ3���.�$�
݇n��T���f4��ɐ��AI˦^>��+��?�n�%	��'DM��!����N�
c��~��\8r�w���������~��~m��T����)w��܊ʄ����@�F�-$Ƌu�8��s���Ҍ|�iKw�qP�-
hG;�JV���SI+nb��&���� �҃�\�׶�U��N6�<�����cR�yy(���T��N;f��yj�u�u"\i/@�EB;ϼ3dpk?������R�'��1v��a6��3�Q�3����#�1p�g`Ǌ,B�D���}lbpa�?��^�m���CtkV"g��*�`XJ"O�9~b��pJX����d�ī�D}��9����[0(h�	�bƧkf�(������h�x��_�S�ܗ����G1'[6��I�M~41y����>����#-��g-A��۱��)�J�"�ߢH�M+Ks($���!��M�vG�Of�G5Z+�v����`�0�٨�Y�W���>�H�����I/�Ln5�����J:��"+��̀�-�D�\�8}	�z����]�xD��D�� ���[D�$���U[iS��nr_e���!!�ީ���A������h	v���X	a�(�E��·��ʅ

p酽A2�R�%�qm<�� Bl>0M�XK�5�aP;?8C�<M���_m��y��^�S�{]�(C�{��y�~��ZS�	y���h��9����n�$]��'K,?[�j!�J�1�pT���1��0���'�>\m�.(�P7N��I�� 6���A��_��}��%	��9dD"I�"�}dp� �AbU�����q��3�Wܙ�>���u١���}Q��Q*�Иt�F`����ܼ�`_ɬ�@Ԕ�m|g����:7�rm���$�t�e�kj1�$�	ق�� �l/���{;9c�Ρ)�����W�G;�qI�Ygzz`��ub!��� ���v�����f%l�HM����gr�(�*��N�ĥ��ٶ�l+Y8�\����x������!�{e�X	��a�r���s���'U��`��hF��V��A�ō�j��9nK��(�W��)��F�BȽ�ܚ��8�r�՝���yFo�w궛�S�l;��we�(��4� �Gەg�vc ���J�	�p\��y6�7CK8�`M�X��ʀz� �S�boת|�>�̫�ISa�z�J��[޻B�U��V��M�-��ӊ�kD��2�|������v�j�����p��R?s������^�[��៲���MH�5����*k�fV�7����z�'|F��7�J`��z�W7��)���)�&,��y�����V`�E����x�,FfD�~��u3����>Km"��T2Y[�f.b�r��k�2m�T��I�,jm��}�J�/��V���/~a��	u���AhՀG�U��Ѿ���pƊ��(d�f�x�}Ԑ�SNο,;Κ@\�ڦ���K&,f a��nŶGap�='��a��c�����r��Dy���1�h�"��y9� ���	I#)��GL���C�����$�r�s�,5���E��S��2ц��e�F��i����O���;+z3�|��W��[�xR�6+�RWn�r��WBI�o�|QƂX����=��p&����]W�~�
lV\6$�:�D�]P=��vKUeP2���Q޵����Q�ç�4tuX����I������Rq�]�'�l�c�t�T�FT$ۢ1���&����l��?V �ݹK��@J�Zw�L��.z mI���hJ���aT:#w�����Q`����:�ɔ̀�_ھ��ZM�J�Хl�d�/��
2[�@$���x��=4(�]}� +$�s�]$����Ph,`9G��&{O�+�AL#��s�a�t'T�B�8)�mm����)�uz�NO5t�xP�I7�r��
�o;� ���s��Ͼiq$�E@���j.X�F�R1�}i
�aq�Z���0ˆ3sE�&lA�CO��.�"8�fv]�7��^�-o���kiQ��E[����'�ܵ�V�r�a��������p��voI�t��ʨ��؀��P����Hq5� �(����"��_?�W��i�t!�g�Օ#wd�v9��@7�q�����~}"J����2�h��xYw�$!mp��mxo=kM��#�3��͗�I/O�Jʥ9���Ǒ�I0a���j@���u}��)_���E��y�d�����U5X�m���K���	4�'��I�t{_o�/�e�ސ�g(����#�F�
O����(f�OFݱ^�i�b|��,�e�$91ԏ|�K��߿/���a%\ ����,����$S$�AV�NP �d��[s�N����۔��E���v�䯮{oÛ̖��#�	�{���ѶTVJ��%p��/�|ԱϞ����:<�
QM����Z�;(�:�v9�]٧�ޣG�B�ձ�+'�����&�O`��M~{qI,O�)���w1��b�wM}c��pK�\�>j��,/W��f_�er.���6]#Xgd�1gF'���uLk B3��k��m�?��a�׶|\�8�Y�q%�g�o�&�q1�]C� C����w�(l���OЌDK���ʧ���[����F�x3S�3���F�+��X0&*:G�`xf툸�_(�c�3�
��{�qz�S9��OoV����w�8{!�p��6 ���샢&�n��n�38�W��<+'Va�/�����cbZlLq�n���d�ZE�f�z
K���ܮ7�r;J����O�r����cҐ�1���ˊ>�o&�b�'th<�x�P�u%���?N���l��G�uO�L�")��gǧ�7Ӵ�v���=Jz0�h�&�\\�#dဓ�?�~C�����׏"h��ʃ���g���l)E��,aZ��E�s�����V���pQ�e��V�o(����۬ǡh[�k��~���Xy ��.�4� ��痊P;�X������q+t�Q�^��~v!��Z�s[�fU.8_L^\��&�/A�:�}3�Dkq7S��ye��D�t��b��[�.��hq`
rɿ��XwÑb�b��a|�u�
�xz���M�ge�iߛPS�:�S���Vñ}4�mqtR���6��(�l��nb�l�g3�E�6fw�����oh���M$��͝�Z�*�	�m�<0�՞H
���ԕK����H���xC��B��=�<-V_�y�T�U���g�/�8l�����Ԝ�
l7tΚ��$j.TT�����CLj��.zv�FJX('�3�M{�0�E�� }���Y��c�7�k��V�q����s�>�������r��so��n�-�N��2D �u�?~{B)1�����(���w�uC ��f�2���h��Q��d���N�.mp���R%Wt'��+Et��,�#%�%̞���	ǔ�Yч�
���`�҉kiL�x�,7��+��U�Y�S��h)eoP��.�M����C�O��J�x�h�����Ƈ�0��{���CV1�18c�Uw>��_���;��<��h����9��R����m��q�d���f�c~]�{���a��=W�6Uo=���W�d�G,��SgN�<軠3	h�7����s"8�_ŵ�){y>��j�;��1�\ֲ ��+6P��j?{J�މ��'go
���"�W�?�I���X]:��(/���2p=��'-�|�E�#�?��K���ᱰ(-�y���~R ��L���~���	�U�����P�)�f�}+Xdcj���2"U�w��EM�'�@?
� �R�z���3 7��pX���0%�pkJb��M�asz�N�]
C�E$�!&4�G�S���%�иXg9�樓� �,ĀAC���N�"�ժc
\�9�J����#-|�b�
泋ȗ�[:c]�q�;��[s�<�������tv�m��Q�����C� �o*����4Z�l�;�I]Qw��w�*U8��s���ab3���i��@9�&��B%���u;j-��P��P(�6�.O� �QsU�����[u��b�x9�y�n #% �$m;GǛ�c� ]}���(���Z�Lk�<6$��4�f
��n�zg�9a��ۻ"���%��E�0��W�3|٣x_湿�b^���LG�Π�!S�!d�rl����4Ul
�3�2�A�r~�mUv���呹N��m!�$�m '����H�Hצ�Nz�m�\}��픿Қ���1d�ڢnL�.�9�Ҥ�#al��Ju�?�k2�����g�E�jc%Bxe>��Q""�?Q�6��a���N7.dZ��R�	��=�^&�,m��a�@O�����T�`!y�l�C*�j��{A���iUb��*��Í�1=�=�iB�?�}���/c�O����)p�j{�$���w�P���x�}�yB�W�K�O���>P>No�KHμY��Z�8:¨`����DO�(�F��\��ȗ�W��6��)_���,�*<�2�U@�ĿP���^6s��8���H��@���4�-�.���fh�����m���C���UE�2�P��ݏ|���3�-�*�Ǫ.�,�v�K]H%���_i�S�v�UYuq�<�:���L�Wә�ژj?&{�Py�����Ҝg�t��Ә���fd��<3���_�oW%��4JD�6��g���nE4Gag�Y3����B�dq�qZ���j8^��?I�����RI�"z�����L�P���b��*��3!"�om��1��Y�4�{�8n����Iw�����b�VU^剔�v�B�g�"��3x)<s���?�#��������y%�艃$ Đ�7/S&<ߙ�:.��:�6����������_���]��e����\�g� ��E�&�-���������uN�+h����(�,�l��A����na�En�Q��K͔�w�����}����p��gT��|gm.bß�����)7{��s=�G���0��ר�G���DD�JN-Ϟ�*=�cR몼ljd���w�	/�`� 9z��|ϝ��� :>�����V(��W��x���j�%	��gό�`fw���+�?B��� �uNy�E��̼+�9ߌ���팓_��{�+!֋I	�m�a�w���������iXJ��r�̀��48^��}v`���T�l饮�+�pb��1~��R���̚7iI�i[���s���D�SƎw�
�-PJ��d���	�J��K' �ݕE�moW(�8���v�Q��	��ԏ����#vV6���T&��b���c��
.�s�]�=a�U/��ކ�W��̇2��*U��v�.�#B�mxe��P蹿�5�9�����Y�W�"�����U���4��U�[��S�}�`����~����<�д�I)��O�& �A��}�/Onsk������ؼ��iS4�I��I����S�*��Ed��$��@�.a�e��;�:&�|!q��7>�H�ߏ�%%�D�`��Y�O5�0�Mv����F\��fiȭZnJ�$��n>�#��U����u�iCb��;�f�yw��QP�/�}��,�sB#4����4�Ҩ��J-���S���Ob�2}�T4�����$�A��:ś��b��n��(,݅%����(ƳfB#��[�[�_n"4���)�G��d�#����<]�χB�M�z7�*��a~����0!�+�3X�}f��ϗ�QS,?�B��-`�b�$M&&����u�L�����o����y78�A��¹<�S���j7C��
, �h�Q�)S�[����6(Vf.��~�/Ux��wM�'�h��t�"(�Nt��Y�~�ʗec�GLI��KU�/qI2�#'2��XZh:�gy(cH=��u������!����i?XuZ{7:o����3G�A��`�c�_��l�xKq��v�<�%�☫8��bo�ϻ�P\����J���m��`��$��CxϨ�6�;���2 S�'�w�{�g��7�F���C�枮z]�w:TfDwE��?�]i!�0Q<'�A�}�OJ��� ׂ���(��h�9v/Al��;n6Dgk=C��!?|�Bt��a�C�%�"Z-��X-�y���x:���u"�<W�<�bZ��5��~�T(3G*.Y���3����$��RKߍ[�5Z�.(�Ʋ�pK�&���ނ��t<_��~<�����	O��$}&l	�G��>��O,���y���B�,k�5w���4�˽X�V6�/�+�F�5�p�N���\�)
��{6�B��y�xQq52(��>-����7�G_�F% ����)8� P?5���&�[#0I64ƼY'�,�p���V�If�Nַd͕0�/8F��2��.lh�Y:�	�s
�Ҁc�u6��_E�gi��7yK��#
��C�h����Zz1=�e JK!;`�1]���+�A����9�����b=f���$e��qOe����]{s�����@V��7� �ƚWI#)e�.Eڃ�Ϝ,�^�M�)�����z���޼�s�N,2 ����oE�'�I;6�3��%�K}�?*'M"���m%)�������{��T�v����e����%]��L�4�|~E2x���L.�b{��
��W:�?��,�n��H�~��.~
�ז�1��&��\If,WNX��+�#� ��֋8�{"徻iK����8����q���ǵi�-ݥ�\j�v���h��	h�؝U���0����DB9����=I�Ր�k���aT�u� �!Ǣ�P�Â�>*�ՙy�Y�2��^.n��Lt;1�(Eg��Z�2��K^�E��D�R��<��<~����H���r��^X"1fQ$�#2��խH�#Mz#�ۤ����SA��M��}#N�-�gO,�vO1y�6Zע��D�@������p��9O@v�e^��`��z���9P˗�w{����.�K��P���?�	b(�����8�����D��FL�Ca��!c�����.%i��g���q�@F���ٺ-�8��tjlT
ӵyG��c�<싰��7�����[�~7v��]�YíZGm��ސgot�V,ʤ�A�0�8wX=�|տ;jl�^��aG�q^�¸�m�<|� ��)�?jС�c�B�<aN�� `}Z}m@�����I�R�n[~F�HCA�f�)�'�/��x�fpy]�(���U̼�g�ه��+�S���;��l�����##�f���5�\KM��Gwlӯ��!
D�B�O�aCq
vؒӈk��A\�L������?� ,RHxl�i�I�mrA��I@��&,|W�~���jPom�W�b�H�Xa��s�A��갺��b%�l��Y����G�u.����)�2�bs��X3�H�eK�����,\���I��㼹p��Î�j/��5c���ɞ�jv&�s҅b[A����h��˞Q_�t6shf���#w�^��M{$���ׂ�1	_eY)�BٿuԮ=�g�*�o�V�Z��5vú`�O�5����S3#�`�V ��J����4��K ���Y��\K|9n	!t��g�
�k��>i}(G�+o�ͪ��+�s��k͐`N�i\�DP���d���E\�.dJ��Ӌ8i���e���aN�%�?����W�A<��`�������?��q�� D?1�z?�;���\5P���wIЕ/u�Ew��e� -�@J�p��1b���*��N�[z�v��:�2i8N!�(Z=ű� B�Fo��	nL�#�e����
<�x�P=�6ST0v��ٜ���şl�ds7�3�>�8*v�����7�<��|;���	�_���u�j�.Z��Z�5rN���?�
��i�W�i���K��qve�q�D�:�S�of�xǟh��=��Wxd�
�p\g��2�E���ۛ64�G"�{'�Cԡ�l��%;ק��p��L�g;��±Y�tq|�맻Mt�rŭ-�)��O��Mג��m��5�ߞ�Q�K��+�6�0�a�u��w���̨�!�cf�E]n!b��W!-�4�(a)ѳ!icߥw}��ꁴ$�ן���A\ �%��:��7d�$��ˌA����N��V���,v�ƴ�-`מ)��>�ީ�`d玨Oj�ۂ�^j��(.�rѽ����l*ü(� x��b �S���o,G֋��s�^Բ���#^/�������i� � 5�U(@Y������M��-N�>���8��7�ƐG�ʃ(`!4�>�����+����׷����̊�*�n�D�,4N//H@�g[s[aK�^/E����C&m�\�_'�)_�IW��|D<�k�ڭi&&9[��d�w�]�M����u'z]Y�'pA���ȷ�G;:�ec�Y��7cN�Cʦ��=��Ƿ,�ɂ��!�!
g�r������w�H�8��q�{S��'�������{Rp^v�{�ҹ�`���WH@���V�߭"���uq?���\ =ۉ���"{�o�ef5FL��dwl�1�_K����ʰ���'<�G��I�B� �w�"�d��s�#������i=����0�$�آ�kkv7����*�-D[p�����97����"���rs}ȵ��!��BY����vʼ�������"W�c ��>2:�@O<��EA==3�Au:���ô�\��6�ʼ��SV��%�: <�îs�8�%�k�?
ߨ4�	�x���ی��H�0�D��Ù�='d" ���6��tB7��6���&��Ω%}�k7.u7k�I���vK(jG`�
��,&�	^$;H����Wֆ�WGga���7�L`<+��X���ᐇ:���������N��Æxw&�V�ubf��s�)�x�i�I��GT�
�;@�y��æ��_�R�z��&����
`��
��I�(=?�z��d}���o|=!� L��{ǃɷ�]`�Jr
l�N$2�e���{�_Í�����9(y��J��x��U��$��Q�WL����(=
�,4ſ���e��#v�c0��[����)�Ll��}���N�_�}O�fs��.na���uW������k*C�&�o�Sޢ'F5C�֜-�r|Vq�b}�5;����B�r�B�C��w�WN�,��܆�ˊn�0
m	���+cم�o��w��;�s�����I�bd���5�7��^.��>]nf�W4�'黎k�L�Z�(�+4����H��gJ��M@��*��$ƫ�A�����]y[�:5pX�Z���>��zh��^l�?�v��K|χG��cJ����]�;ud�(E�uu
��
�	����|�j!�?aV�X���$
�LRBb�"�<��=@yN�0 Kt���Kl���z0��b��EdP��F��"7��Ҿ��Uؓ�t�_�G��L�3��!�ޡ};�gʙ:h�U+`[ek��^�W�̍�7h�i�3�Sػ5������6����[p��*�;i�t��{�&k"��5����Z�LDT����<V:��k�\�ػ��B8�*p�p��b�w������ny�����Ts�p�߮s�tJ�]�=A���w�yr1����`�zai��Ԣ�{R�:�{	�b�ڠ6L����;����&�l�jgƼf[
e�@�e_��gI��f�%a���k?�Sd�xWB%�#�v#o�k�2����MUj����&����8X����4�K�eDy�\m��uм�+z� ��D��I�C���CΊ�7�h�F�N�Ӈи��Ń%�1�����2^'oq$e!��ה�(�|ܖr���V�y�u?}c�n
Zq릓��NlNN)����@&L��������p�oq/�mF�3r9��x]4�����:	��%�X�Vg���낽dFNn���siF�燾(&��l7z6F|�Y6|~Ʃ9���Q��}3Cfd��i6�CYK"�f�f������+��$�,�m=�˷Z�Ԫ�Jq�`OB$�aU���~T%�  ܄�ڝ0)��y��{�w����?Y��b�.
��	IYQi�OB�9���t��
��G}��®J<�?/Q�Z�D^N�@����E$��`��;ݚ�s�K[|�G���j�mEm+u��ç�����S1�)E��,�0���8�q�}.�]��zS��P�h����l��;k:3|����� ��~�hQ�2�$����O�
��R�{�0���zݖ�Hl�����)X��"���掍����hF�d*H�5�>h�**2&���}4�8nC�Q��N�\j��J��N[��o[�}�0�S�j�
Y
S�t����~~惼T�
Éx�^1sWףm���y�$V����>��Pۍr���
h�Y����c�����f!]ot�E�ʸ��{�
����#�~g3�и�X|D�m�Z-���P�kQ�a�_�W_������@uc�7?$��ёJ���������;�"��&��-ϭ=SS��I���YK�ZUo�q�@������8g����x%wn����a������z����Vy�_]4y�k���pp��x�l(�� <~1=����$)|�3��/�t�Qt�=��������_=�p#�����O�©��~O�q����A�D����̧�ǻ���Ka�l���k4:�gS�X�����-�Qw=��-_�;��P���8؝ӣJc�.9�Wz���Ώ�+��_4�H"�J/�Q^܈#Sk`\���鲗�M�9$r�T�[&�eɊ�2=u��0��$�͟��3ա䄝���'R�iC���g݂�9�������&�	Q��{�ryFGN(ɣ�&����~Vs�V��D�Kq���AL\Cͤt텏t4Q^1�C+����]i�H��b�C=ר�����v�����pO���))���2�Zh6Z��9l-/�[B>�F$i���+��g���Ñ� A�w3,�S7����.�wn�8Z�쿤�0��ow��}˺<��[T?���n��a���7�Օ�W$d�����Rz x�!��r��%!힔ͮ�ܟ�:f�J����e�BD���u��Ｔ:uVwM3��;�l�� �1w빛p.��~K��d��E���Y�y�2ߨ�0�cE�O���`<��*���*�w�"��M�SeQ�;���{��'�OY�mb-�C���]�7��[��������n���Q*xd ~IҘ�ź�9<Y���,����]�_4B���q�����ض>"<���=�oJj�6�^�������W�`[bIWb�>���4��1}�X��7a�|��;��'�s�d��������nF&�y�-�(N?H�g����x{��9w�0%�
m.��۳�*�B�2AC��+ܬ���4 �𛯟�����0������v�+Q����-�hB�qgH���i3[�)�|u�,^��o�>Zj����Y̶���أ-O��n��WP�qeSQ�<kWA����X�>b0��J��.vu���~A�G�^��Sˠ�Y"�Z��'�ZF$:���Y�lbדRx�t̲fQ[�$Jq.k�@���LT������)�X��E��1v�V�N�{�h�� ���I�����X�B�l)�:��^6\�ɕ����#b>Q��K�FD�x�����	.B���{,� Z���9���G�I�
����m9�Wiu����D�d~�������g��6���
|-+�)Q;��xk�
�5����<����>Ghmm
zy��6�[qh�]E�3��V+(i��Fz����Ɍ̨$?]c�U�`l[	Ξ>Wx�I�ڥ+W:�RO���������I�9�)w����>�m%\�8�Np��ڄp%.�9t �-��.Ґ" �$��j8�PP��V��q=c�ԉ�.��8c����;�m�n��3S?0��U2N���e%�W}��+��z3�F��b)a�$S�X�VJ@kK@9��R�ɟ2���W��[ScW^)a7��i��Ŋ����{�h�[���7(:�Jc���3'�\��另á��� y�ojQ����`�R�o��Nօ��xɑ�͜�iE����ptr
���ν����{�ȓ[H0��D0�K�����\�f�R׎��fhs+E����a�uUgD�?2)[ g�T�mM�A������'���u�\ ���'��@<	��DI�&��~�����H����<	�����0�Rn�j��;������B	n��R3�����?�5��])8u����xʻН�*Vgs�_0r|��{3�_�$3�$���$/��.
���[��d
�W��%!�)��®�E�v���{Ƚ��Hk'�������٬#S)0bX����|�nj�R$ـ���LM��� �}���8��!���g�޹�&�̒0zP������a���5���̨u!b���;+��+������
�eDde�w`���sGf�V����	-���5q���g��Kq���<��כ��9����ܲLg�-�a'�ߊ$	A�<"���W{�h]�\e�8-֑�q�i�s�������A��$c�Ϳ֠o"3ּ��u^$.�m[D����yK�Q��<��1�<�͜��R[6ڕ�o��[��qw�|��G6�s��F�W��!���U����!��@�i\��a���lׅ�P����p���>�����q3E:d��=��.��.@S�\َZT��������2=���[���\�}�ؾ�
�P�Q�x�	g�ׇ���6]*�}�L��f�`��`����f?��?+D��u2pC]b�uLT.����_�����6oS�f��t欸,M�2NnÁ�k�\�o�<E�?�38�.�^Pp� E�R�t�8Mݚ4���3��	m`��l����O��6��,c�b�ڮ-���-j�А���5��J�s��k�Ŋ�=���kM�/�[�\m������zD��t�G�z8���u�ʵ儹���(�OU'�)N{ �|cM�/BD�E@L���;��j��\��>й�'�~ކ��C�3���	< B�f%�ۦ��Fo :3��g3=m��t\���`ǉ�5��<��s*�?@M��޳�7b�D��)�����I��}�,�������I�R�������}�̨�Z=<�g�`��nO�5��μ/a}��31�.ŏ�K&9��j�����w\��2|BO;��.,�O�����w(����8Rٍ)��?�r�Gg�`&����RG�p�k(b�`��m
Ta�=���uw]���j݇���'��LP `jE��J��ʔ^%�_Ҍ�dب�<�#���(�>�������$��a��U$V��<d��<ՎT�*��b��k�i3˄V�=�Y����]�}�x�rr�b����v�p�Y�Z�%�uY����v��b��7C{�u�_q2�> ��͌!J(����u��iin�II����47�������ƺ�ɰM��KB]x���T��x	({GE���S�l¡��Z�N��5 �(�T���b,����T޲�7b��Ae�4�I�8��hsXN-w�K�<����R���jLT�I��@v�i�3���bs��R��ϼ{�%�g�F�W᪼��9�H�R�Rq�X{Y؈���%j��L�������.�����
7���;t���U<_?�qc.��`Q.�%K�P�0z��-��8�&������B
ԋ�c'�2���o#e4�����*��\כ%3xn�=�@Z$m
��㸄�P�nƊ�>@�\�/�X���l�zb�AT7�qC5Us���,������y>��>~�q0ec�6@]M.�^*�����JI��mF�Qr'���ʡo3�'�#s�ڴq�>�>���f'�?���jx6#�Y�Xx̴xm��B��3� ��9����e^<v��[�T��E���+�P�}�w5��G�|�Jk^	��6���~��{&�R�,Aa0q���9����R���
�U^>�T���!���Nל����,�����= 15��¸�2BO��ly�nIh��6��hv���MS�|����FG������h��W1��;_�0���}[��L��G��д2�wm��;�c��ǖ���{'Q�}N�o0���*�2ח��#Aڤ�k;1�^NPa5gu�\()C�9��s.���\7l�v���
�iO�k�g�����~�H�.��wbjl)8��ፙ��� ��^�\p��yW�Vb��i�g^��9'�Ŗ^�ՔU���U�ފݩ.'(A�>u�_�V��+��L�D�j+�Rߑ����<"D���<�NH0�v)E��BP��w.v�#O.�0=������U��BaR#}�h��#�M�|H���(�v7��#��鑪?��cMOh�i!XlZ}�45 ˴��#�O�~k�|�4įG�s��g�c��M�O�X2ɑ[�O�p�z݅ҹ�HvO��1<D	�T��ː/P1h��?���f%�{��	�W� ��@VZ�������h	FI2U�"�cO�ty9ɲ�qiW�810��l%�X�y������c�2C�ꄪ����2���G��C^�h�>�������xH��Ps?��T���汕Bb;������3-���v�P�����Sx�S�y��dw:}=�A$zhE12'����ɼѕ�I�u,�����B�m`�_e$��YNG1�~l�A��l:����v��wU��I��^���5	,���W �md`�?���p�>3^-����x�z�/F����(�rҙ}Y2��K;I8��H�����EO����.�P0�ȼ�����"�
u��f��ƻ6�\�9,��{9'�
�����D@M��
>1f�U�g2O����<�����켢��F��P#��vEz��_�7:�@[L��c��2DKQ���9o�1�1+<��������;5J�t��).���EZ���
��7>�o�b���P� k04�QP�R�k1��)�QZ�AĽ&�
F `�d��ꅻ8��0 e>�U�������/��
���e�~ tb����!Dh/;QS�}��<�sq��{H�6�D������S��z�.�Ĵޙ!���c�b�9F 7�"�J��&���&��{/����s㎆�`E���AX���c�<�,G�C�o燣x�oF��=	��S���y6P�aAp���^a���gϜ�M�B���D�\3�_���.��)��m����8�ډ SX��w��D��)bCw�A��^����*�'0*�h����OY�bPZ�R�9I�e����#��	�k��a�ٹ?�îq̏���Ӓ�a> �}L JϬ:u9��x�ZM�(�B,<m�3%�Ƌ����O<J\���< ry5`hfV�����1��nh��p���'KǢ�Ux~�_&j�3�a*�i�*6�B�V�!��)-(��g��$�T�Ɛㄅ�'��h�>c
4�ښ`�S}0�,�������5�r�#1���G�h	B��N;~?p6n�v���M�m�T��l]�8�Ƣz���c)�^ҷ)���$�4�c�r����|d���X)@���ߢ]�=6�?9�w@��#�%+"����cb}��
���*�ɹa(�tFG�a䀔�7�Q�v�����	==f?W�:���=�c� G�W�d[�2��K|�w��/�6�6
/��PqlV�
�W�Z;��x�:��y��si�o���])��8�D�`k�Բ���^�N�~=��rtv���6nV-N�c�~9�)B�q��j�NX��3��^��r(��,-�@�Wށprp6n�JU�O0�.Ā��V�3���q� n7<�)��*ݢ0�6����P�Z��Y�n���;N=�z3�1��� �&')�;(]G*�j	���2Y����+?&����wK5%�y�
X�Us
��a��'%�8(���G��&<w_Ic���$W��k���˧��jVp/�r-ߦz@�n����'4z���j(|/e:�H!�q���]�i�w&<���;�OX"H�^=�}deQ2���hE�g���$ ��)A�A����F�o`�?���bC��=��>s^I[3t� /ְ�䠣���-�t�����(O����9�6��B�S�q1���LΑ�_E�m����L�Y��bG��*Y �˧�+D���S�`Uq�_�U�>f��_E3���Yx��h�-&���碦�����}SxAP��YJ��϶����E`��[Y�N�ˆ޷�3��q5wP}�z��N�)��=!���ʶ�f�	��o���s�����S�8�|U� ,�i0��~Q`G�2��F<�÷��B��r^�]>( ��Z�(�����h"�)\�Ո�+,�3yڏd;YI�wgQ[�Q�F�hm3���|/)�� Ӟs���)qk��4b������	����y�{�#v�N��ul��2v��E7�i8c��G	�e�DT��*ќ�$�^�9�D�#!?�M1C���K�vjGCQJ�p0��i���Z��D���b���n+ n��R��J�?dMg�3և��^�K�N?K�%pkt	o��i6Ġ6
.!�5E_��Ј�d;_��3�f��#�ލ��L�-쒝��>�{�^L��n���KS1�~SPe�-�c��i:Ǎ��D�Ij�^�[./aƴQ?�&�wyX�r����e�ԗE��A����t�1��rYwqG�v���N��P.��|T.(��At��&���O�Ɩ4�ֳW;������8�2�����ao��0U��ֹv���_يF���{Xx^�U`�M1�fQUP������M���a%S�Zye�&$e3�*�z�a?�]%�i��4�
�*�y�t�8��m�Gj�V /�c��af�=u0�n�q����YziF����މm�e !
�_rg�7<�~\6��I�B-�AEz~P�4�fY�ar�@����>�i>6��X����_��u�s�$���e>�S*������N�Uw�b
S���i����Òu�\�ո�jb�S��{S��&s�m/D���n�&Xrn��j"�Pq.d��:�r\h��϶��oRMD^l�k���zJ�<n�?Bu�H�}��Q��l2[\�]�EMQ�SzWO�@������o#ZWRI�����QoS�`�X�Ƚ%��X׽�Z}�s�'�Y�U*1jB���*=��>��M��;�WC_o�(��tqQ8��vS)�iud2�0�lWRK�(�i�[��W:��h�� ���2�d�\y�3�x(�A(�؀���U-�&yi���γ�^_�f���d�Ď"�����5�Z\@�XUһN(�w}��a���s��b��}l��J\�c�hAYh���a�\v��~���G	����]�Z9{ae�pqj)���<���;lI��3]�#���a�����B�Nn �q,3%�*��eup�{� i���BM�/��I�����,˻����/.ϻp��+�����L�:�؊�?�ɸ�N4�\�n��E��G�F���z��}�hx�A1kh�7�JS+��X�^�a�R������ਙM��#HZfs�݀`�]�3���J2y�m&��#���x^F����Fbg����w�D��!M�f�ϧ�%a�����a�Hy��;���8b�7��S�&p?Nʗ����Ns>���tm��0*kuRj [�Z�a�=\�04��	2`b��7)^8��}*vD�*t��WE?�=ٜ���rSn�M��RP����@>���E��9;zmZ1�p�K��q0|��GS�C2�'5�-Ȫ]�Rs�S)�l�*T4J�ʅ���cSZ�n�����$�%z���5-De�d�{�p+�~��NJ_����&������)��RWK.�(�y�3qȑ�i~�R���ϧ]�� ��g��ns�k�Y����=�3���3�r�qa��B>�WN��qU-���w6?��_3Ҧ$H'��ImE�u��4�~R�]X�9Fe�%���Y�g<%�������Ə�C%9!K�_��
�m;�I��׼���8��"͟�6���KEim��S��RF�`�e�c���*Ʉ�g*H9S#S��d���r)'5��}�#wC���q_��l��["#���,��
�	�E.��y� ,Tju���7��9����'E�����<���5U:H6��Ѡqx|(�q㧗�q0$H�# )N,S��w��V�ZޅiA�U����ev8݄Гp0tHm����}U���A�b����Ĉ�P����HMG&��zz�
Ⱦ8�
�M	�X�M�Zd��T\y}vH2����[��-I��֣���4��V�Uo���:�����U�c)�SLb�� +�W\A����;L5��s.q�O�
�\�\�lgz�l���S����@���wH��|X!�K੎�o��ѡ��|�s���3�*�w>���Y�P�+ϢA1�'t�D�?a_���{���{�������� �o0Y��s��p�;�U�{H 3!��f�P ��z-��0�}���J��t��a%Ԕ���E��"�x����{��"��D�	��#���`?mr��s��#]?�������2t���i�� �(|Պ�~n����ߐmM1�v��3�q��O��N&&g��d�4���wx,��{�К����PI�n����w�̔�?���g
�f6��i��L�����&`���q��P�T�������R:�L!p���U�u�ˇ��Ο���)!n�*�v�}�yYb����,���!����-#��ߥ/{��G=C�%Z��2D�0]C�Ĉ룑��Z#yF&��BI�(��.mqh�s׹�e3�P�.�O��)��+�\��{w͝L�˴7/���}��;��@R��	���o�`�k���B��%w�E��.|B~��V(:Y��0�Շ�c͖A��Ϊ�	ck뤘�Y6�!��@}	`�|u��Zn�E�"kPi��A��jv��D�B-�<ϘK�����g���ՂԹ]���A#^P��]�w��[�vm��4�we�\PD���
�0
�l�P؃o�f�ڃ�?���k�=�ä��w�#y���-<<c�j*���t��>5�_�s���RʷB�YB�?��c���'�oR��[�����M�t���I�0�bC�_?�� dĿ��m#�;�?)��_3I�0Tq/�e��A$FKԨ�(�KJU� ٦`�r�G�gFH2�tNB�E����7E&,�5�J��l�Ҳ�e��R���Y� +���S�\�P�����A�
^mx�ʝf6ݡr��ȟ;��]�~�vSh4�Yqc�Z�
���'�e��l)����m���
�t�O�+ݖ������DWϒeg��0ȣ��*�/���HP��m�ۿ��@I�t�60�E
�s+������M�}w����	�����s��})<�P��]@G��k}�[M�T���PV:��c��5�[�g��OӨE�!�e��(f'�f���,�)���r銂Ձ��+B�)h��7���n=V�/h�]:�1{���E��}�z�6JA@C��Ȯ ���k+�h�b{��N�ߛ# <���]Qq��s�����.�ek�J���Oy�%r��.Ba#�v:�Huj3Ɛs�&�;���Z��1c�O|�!�7��������sf�օ���T�+*W!���W��q˖��_��5*�V7� )"z{<|����>��N+d�� +��P�ʾ��TIWX� �ۏ����R�&�u1��	%Oꊆ�M���t9��<Xk�5���u�t=��hW1��8���mcu�i�GpǑ�.8��h�I���^���?�G�������Vd���Qx�@"��|Bw���	�%��1��]��A�(O/�i��ͨ�Y��F�]2�f�T�Q�՘#��ѭo�&��@��SW2����XyIz
[՗�)f�I<��㧁	MPy&e'��ө}�
���ڮ�^Q��;�#+t�z�`@���J-���#�̒��T�I��a�����ׄ�k�d��E{�_k��B)����QA�\���JN��+l�\�`�[p��i@��_bQ�#�l�$nۗ�����L��Ec��y1����K^�fB���PJ��&<�;޿`k���������|_�%��B/������|,��ϯ�_�=�H���-!:��"1�[�pBt횶D�{D�V��ER�?QqNҘM�0>�e��{"�w#��Q�_!z�b��5�%��]�0��ߋq���P��i�-���T��V���<>-���5'ux�k�0����iF�"��{�&}����հ+!a�Bf�a�r��BD)�<��5G���V�t��
�KUf�q���O��B�{��.����I��>�� �n3�o��EW}(+��$-mNˈ��"8�!?������Pl��|8O�jyF[t�{{Ǔ>&�8�f=��2 ��ַT����\a.ǒ���q����h��(>9�%���OY}�<nS}V큱��|,���a\$�f%/�[~y��aq@�I����䡡	2����܅k �`{�9<��>ꦝ�ק˲���۩(�Ҹ�VS��͔yqX�)%�T\ pw#�@��n�Q�h��ׂ�@DGU�DN����8������b�Z��v��[I��(dA�Y���M���\���cR�� � ���[Ԣn�1cإ���a�i���Dn.�&��ɏ�s��nšk#s �?g*�Hh�xC��cca�)ů*�*��q�����Fb%a}5��C���,����6���j�ҡm:/�O�
 Z_�%YD���*h�{C�.�t~ݯ�e�r.B���ژz��ߤ����!�{h���_�����S�\^���q�*�-��1�@�D��㲗����IՄ�cpXZ�0<�J�V��o�PQ齁���졪kv�^>���9W����u�kR�=0u̝\��
����ם�leF4�;۩Ds_/�׼dXq_G�ȩ�a��U7��f'�~�����À��N~��zSf�H~��d(�g�3���D��:�AxZ�[xQ���\4�A"�C����)O����+���_%�%DU�V�p!j��+
ɥ ��[�A��^[+��8�D�r��M8ճ�'+-�i#P��y�#��0�ʜ��*A�lJ(B@X���7e��k�o/�tl�3"� �G��!����"b2�5ع��&��A)����m��!|�y�J�� gp�{iu��r��/-qr����{ҬZ��WX�V_X#���;�#�ĶYO�Tޠ�'�!��W,7	��d���?�X".`����푉4IB�4�9%�10��V^�^�[Gu���
u9)r���XZܰkf>�Z��T>�@���l`�k"Xtm�%��*>�2�|V��,���4.�T3�#)xڊ�e��gaÔ
Y�~L4 �p��T��Rx �yi��nѧ�1�kIhi�;�����v��C���ʇ7�88T���?�
w�*����ɗ��@�s�i�� ۪�~��H�c߾��(��@켙&���U�Oƒ=YF�����0НAf����#��4^q��L$��*n�sQl����s���2�?�x�]�����`?��:�Z���@��c����{��x
��-0�V�s��!����D.���OW��������yz�|�*�u+[q�����\�_��� Q�w��Ei7���X�36~>�L���%+8xw������t6y�8�����q�`���}�EE�}�K�"4��:T�I䱶^ ��6�:�>��*��q�)�merՑ�u��V�cRc����U<o�	3��	�H��i���g*�*� �X��y��I�0y���I�%���p�3U1������ĘZ�����y��$��գ���e��S�2�XK�ǻjP����(��?c���~�ǐ��h��s|e�љ��/.(�@�8�P�۩�N����cɀH�2�!5e=��$��^��?��7C��G�- ���<j֠�
���b�C�.˳�C�2j:2��j�T◎�~m�W��v��(���T�i���K�����ˡB��K�������쒁=3X���D���f����E�x���1{y#O� �������x��È#��m��I
{��Wӆ%]�L+�I�v�5���ԕ����vpǄ�̯��t���.S�g^�6�辝p��Ao�ֻKW�)���K "�~��u.��Y<��s��HՍ�4k�B��,��*�8�Y��V.7R)�&�m�3�Պ�b;ތQv��
� x����б��u�L��,	�Ș�Z]��vw���	(ݰ��������SV�v��-�A�U,��&����p��PF F���v�	�}S	�K��#
�F��Jl�U	���T���������J�HU�g���z�^���f�oaƁ_������󒶭�'����刢����U3���=S��#Y���%���S���Uo�t��FR�d�H�U��~�+W��N��SQo��W�~�����"N�Z�Z�HK��A�.�6^�ڛ�9H�M����1"�����!�2l�բQ�����<~-����-t�J\��|�k���1��9��6���#��a��jL��dYdUwK^R��T�8m��J�r��9����DIg�	���_��f �j����̩'}	��Zfệ)��(��ua��'�����F���:�eUt.b�AGu��zw�l��y��6������C�S��0oI	j���i��{�M�Rz�1�&ҭ�$�eg��X��s�!h�|$���,\�u�i�t��i~F���S�>��E�ˆG^�q�a	��I���W�_1��L�yz=�M�.�M6���xà�Mʶ�TK��ۓ������g���ub�2H_����q.�$詧�4��O%>��	:��gCo�5��V.q{PX�σ]�b���(U�t�iQ�
	{a����Ț�K�#Ix�#���3x�j�,� }l1+��}�t.��Kb�ƚ��P.�~�<���\��57����2']NՄ|���8o��g@|��6b�`�0l��ђO����6�M�1��p��=B>��Io���,�"�.�Z}��9��/6m����C
�g�U�A���-P9�.�n�R����'�h�`�"���͙`����'� g�~-]��g�~T�[�b�MhA,���	�~G�σ|���_�cW���
ͪ44�I�@6�r���t�Hoqq�&�f+!�j��c��E+>�f�W��\^ ޕ�`���+�=���ד���
t"��{8�xh��v�*�"G�昲�fbm8�Ĺ�Y��՟�KR {�.��ةr�C1EK��~��C�Ay%�s��S
��G��a��QRF�ޛЙ/|�I��Ui����'D:^���]�rA���8'�!�y��P�k��M|��)�EȈMV��GK�}�-&��_j�h	��������u�5�s�2M�DUX7�J>y;��{��O^������G�_�E��<h��O��	]��\�oXp�d�h��LLa��wJd��ég��t�zY����8ib8['4?ٰ���/��@���/�Q	��e<�q�'Gq���!���m���݈)���ߥK�����+��� 毹O������ޥ#F7"�Ƥ�����0ԗ�ŜGCFhU9���V��Ѣ��&���A�F���f��9â�s��E�#��ǲ������j3��� ��=�}G�AG�CE0c�vź>IWq~��b�}�ޣ�]�'I��{5Z�h��dN�fx�&�[
产��ލ*xP_jA>21X����X�Y�z�H_ln���>4̞ܵQق~}%HKn�r��R}��,�񝾵�$Y��X�)k����:�ݠ�  5��I�$q���#�i��H�r�'Є�snQ	dDBcO0�/��C���is�#��ͥ�����x�T�%�V��t���xKLc�[�F$� ��
���y�D��4�E�yK��w����;�QI>F��b:���f��E��ɔ�ڞﱭ1TC=$T��uc�g
�r�����[�.-]hRTbu�л���6�P~ Isz��ʛ�-�D>�o��P:��b��L���Mm�����(��C�=丽�H���Ȳ���"����$L*�ox�)77pX�|+Cb+�[��%��[y��]����(��-)8ಿHM�h�a�_=ok� �G�o�O3�A���w܂ɱZS�&���8K[&p�5����VmD�Yi0�0C��E�fgI�
ˡ�l�M�p��σ;2_�����D�-��a�g���s��u���ؔ13��^&���+S ay����?������ࡠ��F��D�x���7�@���w���S�G0s�����V���i��%h���-��h�8;��)���޵��4���1�4s�,S�v[����ʙ�DJ�o=S���vS�®W��L/�8*�T��`���h7O�ah�����g�je[����q�ܖ%,��bY�\��3O'D��_�m2�~V��:Ϭ%��G�v;B����Q���v�[y�r�W�"�ni�d�ݼ��T�_%|/��2��hT�����BHX���)8���c�[҉P�Z����:���0���{q��Ř���5��8A5|���݂^Ȍǁ��Z�+�F�}\/�ߢ�>BXy�/�vi�;ޢ���
�6X�/8.���B�e�5&tv/I�N��ƭ �[��OR��?�`r�T(L��C:�@vj|L<ӊw��8��wR������F#AQ����.א">"[c��5�I/���ei0x��0z�L&�Y�޿�'kM�IMf��}�"�ߔ�2?��V7kD����9�Z����L�౩7}T$�d�vg��}�ó�G����
��G��DISy
	�(����ܤPi�n�N���9��y��T�̉" i84�1B��Q��H%W���Y�ko�n<L�i����l�|ۙQ�W�������.P�(ɸ��� ���b
d�]Z�rs`(�3��7��<eWk� �bM�����c
�w*0��=��m�M�3q �t(�A�v�qg�.�;��1J�7#�d:�w�O��8���K�9J�����tkB`���1�Y�/e����wט�;2���)~gw�8�}E>P���'	��̝�"���e����6�'f �ٳ/�"��濚��J�m���<��:�ߣ�%ܚV}���Ӷ�F��r�8�!��Y�[G2GA>��)����d֦�f.O�[�m�2f[s�0�(����Ԙ���(=U��S��4����{�X� uu��s��!s��3�|ꆲ	��'��9��mv.�6ˀ����\��i�ϴ���}�8i��E^�w�ʭ��4S:��up"�]���ج�>,�e�VG�E���	N'���}{Z6QqЄ��C��%`���=���78"=�]�R9}K�q����
j���"?�m׊I/�ʕ�!
#��n?�J����K��B��~Tk���H" ��v7χA<Y�^+t+���cvp�.�E�N�������d��0���B�S��/Z_�uvtm @q��� �9�=�)�9c����QXڧ�)��DFX�i�0�� ?8����ڞk�g��-i9nBz{0\3��C�'k[X��Qu�1�Y|F�h,�`:!z��aף+RU����u���23Kb�	!N5�xc��>K_�I/�}h�{����`���j��/5TM���PM�rtה�]T���#�Ք�W�zi$��N(���Ћ���I=%�9��h�]���_
:x��G��@�ۄ80 �,l�2"�jy���q�HIU������rˈ���w3s�J�~�'�ОhIƤr��e�)]�w����X�W�{6E\Y���6lǶ_C�4��/.� �$I���k,8v�t�P��Q�E\q^��/��ƀ/��
�`�#z���H��sб���醙��g&�hs���3�,��Qp@ �e�@�6l߶��~�ڷ�W[K !�(.�o���;is�Τ�\��� ڝ�������s����)�4�ߞ��NՠD����I�ӤH��,�,��������܀8��DG�mғ]���_ߔ��*Ҟ�	
�+d�hn��B�5c�A{�c���Vv�yC|XD�
�KѬ����Y�0h�'�p�߁�;"t��p%
ꆮ�\j	9ee�#����P�{�$�ksq�H��W��M��!��<�H5�_E�z��WC�Y��.� d��.ݿ"P��0/��ץ�[��UNj��#�A��o�-F؎�P����c�x[�ف�/AQza"gK#�M���s�����_�=*�x��4�y�%����"X� m>n4��B,a��4����7� ����[[3�+��,.�We���Վ;�
�Qv��v��d��ͰS�F1�;eS��Ch4��c���X���D�Ä�0m������
����~�I�t.[�N%�
Z��ND�@x��	)j��V,��?�Y�aS~򐷍@q���b|zIC���ǂ���������1��~���{r}#��Pݣ([�j�����]�<�����zE�w[��9����H��d@��o�|m����l����J.n�NcƘ���f��e'��t���l��3�h�֋���㨚j��X�GT,��CE���C^(���s��i�(�`�ަ�^]�/��oL���)c�4�!�Z(�%����{%�\g����M)�ҿ���uqZ٬A�㓱$6��(Sr����\_^�Y�n��E+�H���#_Ѥ�A/���@fqt?�Ԅ�i2`����r;��D8b�w�(�|bj��&�>�f�O(��=�QWs��^���
y����1q�u�#���N�'��@�R;���h֍��Q=�SZ�a��A��q�4`Ji��W���s���+x���0�NB�@	����*X�'�grM�Ô�)XZ���+>>�
�.�Jj!�i>S�Ѥ�?��l���;g�-b#��F1�9Ip4C?�%)��"z�WG]ͻ&^�eD�-w{l�9��@�S7��s�͓;9Af�(���G�~LZj��eRڊ�ӌ���i!���Yi߈�j��};�ݺ�/��/����������E浃v���,�^����.v���`�}��nia�m��N͔�5zE88�;r�Jv��xΊ��U���� I�6y��Et���U�-�?:�D:��]�T��IZ�:�7b��sR�-�[���S�Wk*VYBC_I���)����j*�~S����4�+�KI[�㙀{��(����[�rg	f��z�oJO:�b�5�e��
���*i��\��ZM7j|�*��L�x���bQ;:� ���I��؛�_���{�b�l#�h��Yj����-U�/I�5�aEm���./�$p��8S��<��6�8��� �9��7�r���+M$����:v��1�9��yK� �W���u�����{��y��M��i���)�H����/�D�d�.l|�؞���Ns	�ry���![� ��%��Xy�=~��ڝ4��7�=���+8��H0*��D�h�� ��c���tn����Y��	�c�@���t��a����Ȩ~=\��L�z�g�N�hÆ��}�7�$��st+�i��n�Zo��v>�`>�Y�=G<���Z���������CS�m����l���0#w&�yҤ��b�Zp�ߒ5���w�si��3Z&\���՞#���h3<�vH��bl�������[�Í�	 ��{�pϋEo��݄k�Y� p��	���#>�-Uos�����pX�P�+��3�jH}ƣ{�̤-���,���Yc=�������Z��y�Si��Ę��>٩�����I��Όl]��q��B�V���;����69��F�%8C���h��6��Vk�ڒ��=�MzP�7����Y����K+�(�7��.��pB'��p��ї���+��"A8�6��(�>ɟE�yh�����P�K^Il-��>�5�Oc�Q�c�������n31@֨>��M�ڍM8|0�z� ɯ�N t`Q3��R��i�����FK;�:��M�Glˌ�Ô�T�oa�I����$C�f��\�s�D�Z����c��43tn�3"�°�|���p���+�C\�g!w�6nrnp���Q��$]O�f�B��k���ⅽ�*�6Bx�dP���b,f�&���H*Z�η"��#m�Z�0Ů�yl��^zȹ����@� 0�㽑���QՌ��x�d63�u}!u*��d�"��:��r>�*(��A|n
����?��	��7 � �H�����Ï��\c3��W����DN6�-�~ᤨ У�n�۫�>9cw���`�����YM�Z)^�3VlX�&�vpsIGP���m�F/��`z�3d%ζ����gz�-k-U>�TQ�����3V #����f����`%�npm�=-��(������/���� ��v88�iA7���P�l���	�xΫq�������4fv%2\_���mK����~Gg˯��$~3�I���5$��̈́�W������J�
B����Y��s��a/4�R�8��{.Nzo4Qn�j���F�MW�OCW�h��0Қ�	���";�@�zE�=���+#�F�ل������k�I�3����YW_̖���xy����k����������um]U�~�3=���͜�'��A�D������>��S ݒR*�	��=o�(�Yg�ށ:�*%@���G(�c9,��y�Z�{��O�(i�\L;R��CZ������;N�w9#8ڧ�����XB�)�������B�y솟=����d�����$�H��M�0�Z!n~���n���?O�����������2�Nl�b�A�p�U�j���i͊Ø�ek\׷�q��0�fAHPƨ*����%�ջ�e�G���A�2���{��yuf~�y>���L���ρC�ݝRk�.BF�-�Y�M�iXqc����:��I	�2
�L?q�6[S,	��*��BfL�Y ��"�
=��9}�:��N$��/���ݭZUS�%���:���»�g���^ْ��ب�pv�WT~�)��%lg| Qpq�%�+(/�0�yrȰ5�B�lw\��Llyǘş ��j�8�T��a/?����))4��*U0��F"U�����k��^�`я"��LQ�W�KNL���/����:K�+�3@�-i�ʚ�y��r�~Oܭ�'�m���ID���Q���u��\�tT��4�����D1*�i�3��S����B����C���"����b��*p��	�q���m�S	49N���ufo8)���滫$��~��0��' �(�Yc,����Gr�p<�>E��OF�8�Gf�A���f�wf%*�Geg�Ar�QL����!ߤ�!TϙaF3|1�ߗ�E��@�ay1<3處R��`����SjU80ɶߏ�-˼�W�(&n��X(�7��#L��r���z�1a�z"��)�'�E�^!��#�8�z�:Y�1���)�i��>Z n�+�Jn�ŶO�A={�[0�l�5����iF����݃��6}3��Zc�J/^"G�vV	W��xq�X_��A�a�bƭ��f�q}Cb;�d�]>�3����)hd.��%��]��:j✙N�%Ι�\�130�ú�K;�j�ğP�G�b)R��}�2����4��� ���l���P��*o9�!��]��+ģ�52z�:C����H���ڥ�����5�������QC+��c�F����Q6Ӫ���S��Ms���uYV���)�#�#��O>U�I&� Q'�{)�l�Ϟ�S�������h|�^
�L�V+u�3�)�6g޴�nExE����M�%92�rWƐ��Լ�������y�����f宖J���M���ֻ�y�:<.x�} �����x��]�f�yx��yN�e�WR�.)I����>���Z|+N	�qB␗l.������A��"A���d���ܩ#������o� H�@Sz"�>
L���I��"(>�ZbR6�Q�g��.{a����r���A��\G.�P_ȅ?+ې�qa���ʡ~�Q����c�ݽf�fu����~�������<�Q�قZ�2"��<h�l-]<}BK�eٔ���\h�|�T�L7mm�<f�q�-��~C��٤)SY	@��'o?���m�oeNf�k�q��?=��nZF�S�z����B5i�U���mRs/���CV�m�_�9�νO��h-���p�
����>�+x�i�ֱ1��Æ.K��٨Q�eJN������:��\4G�ʴ�Ms1Z�sd��SF���Zk6�){�h�j2WP����M�"�>�j>�̐J|�, �SU��_�3h�f��G�H���\U��[�����Z��Ge���
M�Ǯo	iu��3�y ��q����u�(�����b�\
����	�S��|�<���k�_����M���˖*�4#@v|�mo߭+!���~�fi��7����V��d�s\��j�'Q�I�5����I��nZ1H��>����$�Ox+��������� ���FK���-��������I�A�YX���".�	|H��WA=�r[�+X�B��O0��(��W"��1"�ܦ¸25Y�;��;:-'�(������h�P�[����!�4J�ɘp�l&�l�o�]�'w)��t�����fT��kꛞ"��h(�H���͓1e�~�4HL�a F���Zm���/g��9�!J�ll�-0�#��C���N7�g���m�7-�ީV�+�Q����i�U�nW�|y\$`��12��5Q@.�G���E���SqDFxR�R !d��,�X��FP~�KE��Ԡ��r9�'g�(!����C�)㹺�����*#>�S�,�p�tbR��.�hAG&3���ֵ�3H_������cO����C���
����r��5%IM�{q�G�ѺV�F3 ���*�#���?c+&L��=�Ȕ�^dI" >�Q���A4�(��m�P��m��1����� ����-���e�d�$��ׄW!���LjE �#���V�_�)M��V��yE����H�bF�T`0.�?�e@,Q1	9�}�R� ��)�Mb��K�n�����nY2G����@Ah�d��۷�O��S�mz�1f�b��-�<�2� 
r���j��'�w���n�683Ɋ�uFk��jo��: ���* ��ݑ�&�"|띾;)�HHwc��$�R.��9'����Ǧc�����߂����D��{'`]����,Dv�F�mBi���v"�9����ZGf�,�
- 5�ky��(gn�Ԝz���C_���e4+cr�W�QR<�p�o��7�\��$�͠�y�����vC���ڼ� L��#Al'�z~���;v�dBâ�t���ϯ`T� .6���#�B��
��.9�1��~��m��em�ÃM���Ҫ����]�w�w��r%j�����j�hƖ�;���A)m7��Y�'�D*\�d{^|DO���432���׺��SeD�7���y�`g�c����XT0�}%���u�by��>e�j����P@�)�'Ē�+���4|c��j[N�퀋��:���"*���-���G�������Ais�fG7#�[6WW'��`y�0 �c�!V@ӹa�	�����3O��&
%�e�q�0���ou��oY�8����~m��W�8m� �W ���[�9��09�	0ݼt�kr�#��G�=�ix��ڇ[�d��ۊ���R���6:�^~oY�v�^�	��AHz�H�@_$�r����l����U$����H����t�}�X����i�cM:�v����V��̈́B� �&~q�;��H/�fP���}_�V��t�13Y�/�:7���C�s�t�]
��v�@g�&�1��':�Z��m�_��<n&)�?��r����CR�K=�r��U� a>�ӌ:��%���òH� 4I���Y���bF�S���0"
�g�Ysb�q��N�:{ڸ�`�����ƌ��od6kQ)�����~g�*���-�zϺ'l`6+����;��?&��K�w�[s!�|2x/m�1�ڄ;�# �{��ʼe`.͖��nWG�f�M�&��]�W"�B`�_�<;]�F�Sh�N�һ��F�D�^��~<Pւ���j�!����=9B����'����*� ��H
�׿�,�*j�9�º^�#��_] p�q5rz���:��[eǄS \,�ƪ�W����L��HN�پ��{^���:/�J#o�N��A�N+�]̈́J�X����O@�QJ%N\v!ǜ��������'[ȹ����Oݳ~A����J�*E{3�z�
Z|�U��><c � S��{��L1��'8���`�A��e��z�(z��I����!7e2�f�Q�*b��sͪ����Tn�`���gǱ�)����_nS�bcSh&�+�?��F�e�"\7����8�eY���>��&9=��+�S����a�S�Y�=Rc�Q�<,��QZ�X�0�C���QK��ʓ|��`�҅	�M����y9hj(\;,'�Q�2�/����8V? �_���v˕c'Q�Dd�"_ĳyݶ�2��ȿj%h���QV��G>G��A��Uo�Ua,Qei�*M6�ۮ�mG��wx�ҵ's�2ko�R"�Y�<e��v-p���W����@�u�L�-���~�6>�g���XiQ���c�O���l�jV �Pu��b_˸���D��>cEϝ%I
�N�Ya���M��hn�	����Y��d�xp��0�.��e�Z[b(!��lZ�s$߃��⅘}?�$	����3Z[]�|U��z�ҫJ�KE�ϴl[�p�-Sc:�*~i���٠�O�W�����n�T�zG��䠔�r����UR� �f�'&0.��d���Hj4����ƀF���<uFJaz�E��}WB8� ϸ�k�@�>p�__��m��<�[�OU-g�o5Q�K9�ڦߖ���0V���\����`�{	��:P^��v(�&�"6@_b��nO�ƻ'��
�Â��{���G��W:���fSp�{^N�n���u5f�Q���vJ�f�A�O[�9�{��q�<���Lw���[�$�1�/���e��6?_ԇ6$1�*8���M���^�9~����7�2R�x&2� �JW=�8��Hy�\����	�z�B*s�Qx�"�O�V�ɼ�F?:�"�D����#"N���w¢�r�nln|�	�m���'x?���.�A2L;}0�G^�� Q�@�iXW$��sh�fPA�_U��.lw1�L��<��L���A��z���;�Ns�+q��3��O�7��E�#��~_��*����x��tJ��^�[u/��A�,�����Bvvǂ����py�0����/�&��\͉�6-�Gg>�p�$��&�񫰏����uw�����v�~$'}��"k$5*X8Y\��ipw�"�W�CB�u��R��ޫ_�?��^�a�����Ŀѳy����V_�Pژn�v�M��3�R����Z7IFIʙr}$�lF����*it��
I�b	�r=���^c�S߰@c�� o��Ǎ��K4�9��M{�X,=�6CX��T��to�ّi����zǳ|\o�<����J]ʰ�$^R�-�X=�Be����5_Ķ^���W?8�C�m1�￬|�m�OTZƀ9��t>�Ci��wT����^vJ�}ˆ xBeǐ`��8[�r^�'G�Ɩ��c��#�f�t0n���m�UK�~�����yi9*%��M|U|���{�>]�!H�VNoHZ-�"Yw���j �P_y��AN�B�)��(��?UO�S�[�����X�+g�ޜ �P�ܗhϧ�v��3�����l��S���trwaRCf�g�=3�� ��<��X���V ��5I}�����  c�Dd�����)�v����faĉ�:a���g�	�:�ճ�|��R���4 Jl8��o�z�@,%�@����u� �jBY��F�����5j��	H�ч���?(��%���lc��u�X<T�pEC��
��']���WZ����ɪ��f��ѷB�������<�2uS�%�̬}LF�;�i�G��\��I8+Y�fQ���6�\ŋ\;B_���)����hh$9�Y�F�����!���BPe��&�9��J�j#���|����C;�}�7�i�������_��<���(^��Tg��v_P��u5�Qz�����:��P�^������%;v>�Fb�VR|�U�Չe"��m�f�Q���É5�h��fĻI[3OI�wgnIֲ�r�"L����"�ċt��һ	���ǈH����}��^�I�|B ��fQX��Q:zͻ7��6����n(�P��4�dm�����<��v^�r��·"GN4'��IW�O� "=�CV�sr�,d�=hhK��s�?��.|�5�"
�l�ˬ��f0W��Ih�,������w�Ժ6+�5�������;Z:A赓���!~(Hm�TG�0Jm�m��\+Ᶎ�m\�6�vg�(��=^�� ��b���w���o�ٟ!v��A�W��\3�D\ש�?��.�)����q#��b_�P$�����W��$�\:%�)}U�R�f�_�n��~����/�h����a���{�ĥ��SVz̳dV���'��1�sb��풅0�����.hC74�T7���~�4�Ԩ��{����wλ�'����j�K̲,c4B�Dt���2��ž�����e�}s���P������|�R����Q�N&���&AU�Ux*�3�=)G4�6�%E|�y��LT�o##�)Ju)?O�T�sI�4�N!�I0��t�� x"n)�� �k� ��9��70@$��`�ʚ����@�S������]��V'D���e������f ���YfW�<���U�1nL$G&1��N�r;Q�1�]�)Occ)��S-���B=���Q���6P�+��)MG�q�b�s}��C_����ަ|S�?��s�(���~��îE���N�ld�*8ץ���]���2�9ڐH�
mvc�Z9GQ��4S(+oW����t���Y�!`�3��5x����
�=ib�����7i#J�|1�!�DM��.�\�+5�C��wq�dNG�Yn�/6��X��^s��J�n�Ll�n+�:5��Lr���;L0�yK7����R�^Ց_�*̉rj��9]��.{������Ib�!~��]m��f�V�u۬ͅ�15�%U�P��;=��ވ�Ͼ��g�/��GUmي }�W򧑌 �핇d��߀��V������1$2�!��x���6���hD�EG�%:����3fN�q�V�QX��k�B=³���w)�ٰ�s����%1E���<�ҲQ�����Iɻ�@�>�4���G�������<���]+1ҟ���pΠ���m=��J?�N��V�[������c�^�K���x����+=u�}rTa+u��Կ%�I��d����?u�73Y�h�Utl)��3��7�пq�6C9���7]r&(#s�9w�3��@�q��/L1�H2��]Uw~���������-S	�T�Y��]L���<v����fK�"�nd�dJ�)��-�K��T�Ԓ��T��%�3)5G� l��.�Q���6[�$�����x��E@���s�����|�7@�L�G��A��5��8\��/a����
|$���k]/\$�/+��]��'41'���B!��xV��.ހ����j��K�x��_�M>ة0��wM,,��W�m���uN'{ 8e��q{,�{}��U�#�'o�����PL�
�P�&dG"R@P9���� M{�ri�J�YX�4Z���n�,�W�y1d��׍���̴�4� $-�y-��`/ș0QV J	��6��(�X��+���(�	���!�k/B�5Ͻ��?(��ze�l�����j�u:��~E����U��R�S^��Us�VrQ�®��cJ��&�8ᤨtD�s�aV<&�Q`a�Q_�y������i���<��[����pZ^�p�ȒN��@#
Л���>�<ѓ����7��v�'��2����iC}0�)5�c�Dh [����s�#%�����uROˣ-�O��(#B]Mx��OlWJ����Q�w�_J��Lu��,�g�4W�L���qnu<�sʬϣ�M��17�qouP���#t׻�m8�~���C��8�\�������I�QGT�	���������m�K���|�U^x��,�q�M�*
��AK+|e`�A#�QkG~
�QCQ���,�P2�:��U�5JȃU�s3���<�	Ԫ;8Y�l*aS��[�`�'��i�ȍsˇ�$ �L0���7�}��Mt��GL��v�"ojJ��PHT8�~U�L��q��6QN�W�#�\psj�$퀂s*�)S�肟ywoi�fe��U
�HN�H����)⾀��1�p��&�eT��d2Q�t���FCV8�B����i��12�q�z�3� 4Yd&���:u.�����χ�x�b���h5ĢSf��$��Db���*ej��6zH*������T�wowpN������
?��='Y�e��'{��i�3Mw�,OdN�0g��1dG�]Ʒ����W�_���4L��Tk|��U?ju\��H�N��E��50�
��M�n���%!�z8�@1�"VL3��2��7�J�� ���v]����]u� �lVB4��~*�Q!$���0Y��P�@4������P��}�`&�d%i|����=�ZV��s@PS�(	L��YZR�ǣ1��
G\�N�)�s!��)��|���ao.��2�1��30��2�D�J�={2�Y.�P�(�ϗH�~��]���mڜa-� ���,/�fYP$��!��������.��pG|6�H֦ma��	&ÔX[��wߧ�{�fQ�	��}�0Cy�C�e}�N����rܘr���y�z��#����A��&�Z��أ�9�$�e2΄C��:���`��D5[�Z�,�{$�ћA��C�凤W�t�I�mW�d<3N����1��'�)��:O��.�W��r7�� uV�q��|��˄�:A.��=Eq�%�X���!��ռy���J�%1 �	���y3F�R$$�.S@��_{3��]�� ��ne��J� a�E1���ʮm�����_�5�\~�WA��������c!m�t��MN����Y��PVm�3��+��� �1���V,^3,
р�y8��A�d��b��(#�2ֿ+ g(��G�K�Cv;` :	��fCWւ��oq�h�Vo�r�͊N��.����<��Ӿ�s��l�]�Ռa�ܢ��˳�u�n�8>)Fnmւ�J �m,7gj.ًA�q@&5�ֺ|��"7ئ�;<�w�A�:
6���$�\:-O�N�AS���t(���,d�ʮ�ˢv���2���f��N]ϔ�+y��O(�Ȋ��<'(�5�1��*gkĝ�G��{r5�@XTt��r�k��ib\�8ቒJH��jCv�eE�zޟƹ��;��N����C#WfMi@1%�<5��+��Y(L�@;�{�J�[J,0pgъ�p=�����2z��.#��ll���WpbG>jB�]��*v������������<U�x�����B���փ[ �.����?ñi��Qv	9��f����T�䰥�	��m�D.pat4rp��� m������`���@�g2�6b�"n!
o�{�v�����q��;��b�u��x0ϥ�mK�T!n�^u�km<M,k-&d9��"�>��įz!��ݾ��^�2�~NK��-��s�`�x�{��1�J�KY����K�]�28*ث��.jP��?����lzWkz�52"FȡM���S�i���+��lV�e���<�܂���X�O�2W��������	�!N�pc���<�� ��P�cGܻd�yu����ApcS��^�Y��Qeӏ�HxrZ���]��r����F��d��iQ1z�^n�j�x��Q���oDʣ�p!�'AaI*L��2[�}�(��0�Q7��nO���L��W�Г 1�x�=��z{=���⤅����}���R7DM�0}�M�))Nl��(�sV���NPu�"��m8o���?п�
*Z��RIN�ʩV^���h:oT䖃u�j�� �����С��ɤ�~�O����+��e;�����y���<�I>}��~�)v��q��O|�u׼��9.�3$��\:�אq8��6�!�#}�Jb0r�񍺪M�,���2��Hs��f�$�F_�D����#vϿ	��j���9ӵ�2�D#���C����~T�D��E
Р�Y+a��4 ������y��p(�t,b&��^~1�%�t?�eb�y~�]@1P��f�M0��z���aFDw���'�����6qk�_1ez��@B�@�_�T��d��}N�� _�@=	��k*�y@�&C^R-Ĥ@�Ѯ��X�F�2-�v��x��L��j��p���ê�gxD+�+ ?SvF�on��u^>��<�kf��/V����<��T?P]�N��+%`V�'뺭q�����u�� S$;�M-��o�N^�ǭ��1&��M�	xbs����"�;��k�Ŕ��e /�Y8�/�jI�`2��p�5���@�<JG�Y��@�R}��_ ����-e'���ñ,�m"�܅&a�[�t���A6��D���,�GS��\�[3�`?���U����:R��8�.�u_�˦�z؛O�6r~�M:�#�3��f�3�h]� �[����,��r�T��HQ��}���ʭX�i�)lzo]-��J	4����"�>�R��:J�"E�n���{`�ɿa.�y�R�I� M�Z����9�����2{Z��O2g\a0u�f*$28���C�s��~U�-�iO��`>=(�jy�O9:�Bډڬ]u�Yׯ��O�E16��E��Za��>���_j%A�4�AM��;y�@ǝ1�������E�q�fܹ�:#T�Ќ��D ���F�
�lQ[,������[w��|�u]�Ts�K��ٳ�����3�U%��b'���'�r��s(w��Gͨ��S3ӟ�����Q���^3�6����3<�?x�a���9�~p��~��؜~旚���˃:Lk�9?�]�^K=�/�,o���@9`�j�V��v��_~������\m����x�:ƪ"/�x�Yhol=d��ɬz8:\��[�g�������c4rh��@z/�*��T��
���'4��*��'���aW�$K��@�3�v�*�Jy�4��k�P�@�Z��#>v����)˿������v���Pu��2�neԯ�B��D���崻kv0o�K���|e��^�Hˉd*���%d���D<L�\�)>W�c;Q[��p`Ä3ԉ�GUR�^���
[�� '~�G�J9��0�M�n`�p��m� ҈qFH�t4�T�P)��4�	#��m�6nb�Z�W�JGС��O��lO
��e�
h_���@�80M�f&s���..��T3��	��f�*�~��\�#����1	�&
�R Fk���ז�A�����Z�巾���JN溮�H� |��c�d!cv-L`Vj�v�%��c?Oȡ�=?�~چs\�Y����O��͜{&H��jL�X����@>w\*#�c�s�jt�u�����7��.P�rK���z5?:�!���0;&�-H�+���sy������`�WҒr��W�%z���A�����<^���Pg��5�S2Vg�O�������k$+i�S�iЋ����mI�ued<�L��M�zUJ�2���9f�6�-R��S8�O�h�k�;���Q���C��$7\�;�FѮ7a,8Ǥ��J�L� ��ÉlC�W��m�
��K޲E�i��J:n14��F9��	M�61��@�t+,#�D��s]u]kD7�*�9�m�H�YHt�����i����;��<U�^��e�a�`���F�(�%9���ă>;*��9�Z�wM�.�_��{�O;�y %)��˼6��	��g��_����j�lK��SH�g4zҠ�=�^�C�A��<a�����-���n~�����?�o�/���"��Qґl�<��DEƹG�j}��ʁ����ᬘ����-�l�F��:��"��QX��{�j�`M����+�-����.*Q�?�*�!H2q( ��0$	q���z9#��x��5G�P��[{�?��\�Q-���(й�W�}�\{ش�⨉g�QHCl�Eۍ�p5){�Z ��Q�wj��t�ؘ�����dT��;�C��ߚ�&@��K�r/|����:�!��7]�U�[� U��_�,ݻ��*C���a������	t� pD��ԁ�?EƝ�䅦Of��	��0�\�ɑ����1!-�H�dP!;h���@�����@���Ф2��}]�ч��0q���c�"e��s�o"��B��"�U99�V脭� S�m�( ����>)��5�m͏'ӏ��BN���2k�J�%3�Y����O y�<��'�R렚c?�SzkߡI%^�NW��ĤP�M��3$�H�e��?߄��bh1����"�*iޟ�d�2P�U��|��
�E�Y�{`�uLH�sX/��X�d���l܍�E�MEO�0�01i�T��?�Eo�R�t7�@�p5d�AG���|9O���bm��>6'?�dv~�^GU�{����	�4���=�EC�P:�A�B6a�L@���-�.N��?��~ǧZ��
f�9���p�.��u�u�os��u���]��c2�婊_Y�)(��0/�ڍh|>W�T� ��ڪ
J�|�\n�kR��Ȃ�Ƣ�G�.�W��Q\>���E��!�֒�?�n�u�������Ai�<�,iّ�@)�S�]<:C���, ϯ޴��	2({�'5�֘d��;eV��j>�̒@�y��!N(D�i���!��>�u	���� l�Û�8%��'��n�hKF�m��ʹm�̐���a�K�(�b,/M)��{N��T�M�cѨb�Zk�p�Ú0 wq'�FaP�%[�yo�-nJ��;V�;�{�����a���m�R��.��pJ~�+�G ¼�f��������lV��͠s��ng�̮��e�j���V�U�3��S�`I�$'�M7�AS���Җ�������ez�	����[e,�*��ǒ���M��v����&�(��C�&�'؜��Ż^� �0���+�v�4�X�Ė �gr�G�o�%^����l�]�/#o�eXT7z�4ɿ{��u�������r.x�(M���� L�qf�:�V�rK�������%����nD�QĂp�ӏM<YMl�PAZ�Gj�`�Z�����Q��?�{Tռ�u�I0Z�	��l�VrX8�%�I�v��9o����LS��R����]�
vrȖ�wC��۟A'�z�؏ڪ�}��u<Ԫ���M~N���CB�����W��ٳ�t�r��5">Bv�S� �H��_��w��Uj�M`��ң9���C H��P��*�Z��#o�rV��a|�N���nq�R�,{?s�%
W%N!���%߰%)�9ARH]]��Y�n�;�U��I'�{��y�|NT�;.?LKe&fz߫+EK�5������ɳ�Mx(�2�K)��N���%K�&��|�qW��N���@T	^擎钲Q�z+�۶��ę�A0+`R�� �O&l�6�'� |A[#�BM6ń�`�]���DXJ�E= �� B7W����J%���p��Qi������x�ß���n^�Y�	�w��2���	(�g&�U`WT�[�t}��b�C�d���M7�+�r�w�@:�b
r"EJ��l\����f�|��$� T���X :o�!^mC��5�۳����"6b=-�O����ܖ�3}ӲY p��Q?`t#�ϟ�2��ʧ�we�$�_t��J\�䈔e՞��N|oFMiWb�������O�ԚC�&��]�w]��즌Z�:�s'd������G�o�cn_��w"��4���|��b�{1�pRW������W{��ġѰr��Vfh�F[�J���M�,'w"S�}]|c,����?��щ����/�!Y���S-�G9�t �kn�OI-�.<|IC.Y����g~R5�R�Ȟ��n���q<O0`$���!+����gZ��A�ī��?���^�A	;�7�N�h��4Z���p�D�YŢz���Ni�ˈ.Fܸ,�~|϶c��ɏ��e��O����!P-�g�v���0/ێ/����H�j�$���ŸMHT����U�>�{��d��!�sxH�mS�/C���
%3Q������7���q(2�섻"�Dކ�<�lu�$۩w�s^!��ל��ȿ?_����q�	R>�v�TI�Z�f1W�S���@�o�Ӑã%�Re��z�ݍ�v!�{��������}�L���c��1�$���ma��X��HL�@e-�u]}���s6.�;<�� ���=��c֜ŏ��tI㪣�{��B�n�2@P<���߼d�ER�5R~�K1c�IJ��է0Do�#&��(5��'E@m��-����@ĝb>�yr H#��9a�]6�|��l0�K.>v���wѼl~�s>���*���v�M]��m�7�EwY�y΢���K�l�;���N��`���hʄST��e�oZ=Ls�C/���f�d��٭U�7��Ѳ��j0y�?���:nQ�����Mu�#�"�ꉼ�Є ͧ��"�4�e	���'M�H&e�?�z/Y ��'7��::Ĉ/����U�䁋������N�s��,l��ճ�w*L�)ҋ�<���m�u��T^�y/:�ԓ����(���n�s��T���ik���^n�#���uٕ�:\C-�Z��KZ�9�$��G0��$�et��Er��޴��i{-��Ddx�Ǒ^8�"�i6��P��ڂ.�쁞���|2%��ٵM���q�˥]��o;�׹a��)7t�IG�yN�@��b�����6���=�#Q����8UK0��V/:��"��m�DJ�#g^!�W���-HMnU�6z��:���)e0.:z#}�Rֶ��X~SX�;��v��	���Ծh~�Z%�Ӈ
>�Ȏ>go����[Jˮ��{��Vv�,���θ�I�5M� �b��J�h���ϝ�j�[����Y����6,�38{��c�x{���z~�-��֛h���"
]7��ت�H1ߺd%;�M{}�� /N��-�<s���O�H���^��F���V�A��,�0�}�W�2?���4ނ �9��>�@_5E���DÓ#ftNW6P�."�j$��޾�/��}�呂udSH]RuO����F=�d��)�� ��dR�74����L�1bB`��!:�X�����%���m�i7�;�<������h���M����Y��غa��&�؉����p=ѹ�1�C����{/W��?,-41ʂ&;<x
-|	����嗖7�~3����F8��i���t�SA샣Tc���%��g��_cuA�aG1a��=X�V>)���Q���D�@� ����'���B��eW���2}_~� r�(*e�zsp�W�o� �p�2T��	*��-��¹�e�rh6���t�X�l�hĦ�v�pC�b�	u��)�'��c��X�7J�P�Q�Ġ��t&�)�q]�SYݬ��3hT��@4p���{��4A�pP0��֐�3��U5)m��+��3����%�~kz��Zt�`�;�r+�d|/l;Iqhj�nR
v�5;~���4e혉K����N����g��ŷ���f��|9�}�x�Eg#m(p���A�MZ/�@���{u˼h��12/.h�.��Y<��Q�j3h~�%��-�K Z7��A�!��;]�V�4*����K��h��m!-A�+�AߖcEmm/��-�-�=�Wg�O{z��"�\�&$pYl�\��t3w�G�,��T;��y�bր�]�ҘP6����0���u[�st�=/�抺�x�.A�N޷N)��Z�8J-"ds�6��'� O �� �d|ߜV�#$qm9���i���ْ���X�5`Ra�qc����ؗ�����Y�����q�9�uT-9���t�i^�a�%����9��V���_h*X�V=�MA��_���$ԋ���<��_�ʨ�Ы����'먫����=K�I��u� ������º�S�I�z
qt��!h��S��!��t�x&x� qs�(�IiN�|�2g���|Eh����>�^cR�Y���I4U�0�� QC�Z��zq�"ŷv��\DОM���W.+�~y㽳L��ʳ�@��M�$.���@�d�����;���'I;O�ں�Z���Ux��./��T.%Q�|6!�1yU�)��D���4J�ޓ�g��&:�E�c���$���HÅ�;�_���Hf�K��Ɗ4��<��܍�|�#4���H�n��~6����He�:�����?��cZˆn_E,AZ^h���x�"cU��c4�@��M8�6u_/�s
Wl����1Ȧ���n1B��*~<��0������NKQh0�e���Cx��R�? B��c}��)�1���>d�p�Ց��m�v�Y_Nl�����l���/�� ���>PP+B�@DZ�^��7���%��2��H�
d��U�ifA�&;�閏������`�f�'�#�~�wԂ��1�cY���چe(U��b�z�Ow3�#+��M �L���
�C�����$[�)D����m��f�Jl9L��t�!��(]��}K����'A�7B��R���Ը�.�fe��D�	&Y4]iyPdd�-D�\�a����|0	�I�$���hn\����+��|�@S+j�ܭ��^���,%�:��Ŀġq3-\��rEh��/���\�Z�Dé�S���	�c�Ie��M\���u��#���M�X�I�4�ߧPn�e�v�&�M��5�<d�ufE��u<q�|;I�����K�dF%Pm����q;�b�hF�<��z8򃎾HkI {_u*I=�.� ��҇�KT.�r�Tʹ��h����Q[GE6�[Kg8�@�|������P�C���n̟��Vy���T y*3ѻ�rBz���xn�S�{��҅�5r��׹��]��H@�B��j���~i����Xp��k��7vh;7EQ���>̉�Y\4]S0 =�Mpa��o����#�Wð����'���OX��O��<��e�;�+5��y�D-��� ?!���� !�W�m�w��Xg�|/{kD%�>�D�#T��O�B��I�Qz �I�mJ��:��j��O��z�*���9�b;�
���화g����,9����JWDSo<[���7oLx�(m�٠gB#�"i�p:1��F����`�ϛ���,)·��ϧ��n\!]��d�r�h�4An\��y��>�$�T����`kH�z�����t�RCc�[�,t��<�c��� ������_��ñ��硚 {gq�|xщA[�� �G|_ژo��/AD|: �B��j�U	Zb�W$ѕ�B�k���݋ėmz��9Apж��Rl�!X��?lI��\�f�I|J�.�Ks��v��^�:���\���NQ��ߟ����x��$���+$i��b���u1.��i��i��t;��j�Yn}:n[���`Q��_G��]&ό	��;7cl���'�肧6�4�3�<ƞ	5��BٲVp�abtW&�<%�����à�ۆ��U�Y�O����g@�C���K�~�����Tc���-��t���Q5U���>`H�*������	S�t_��K��+�kiL:�Y��e���G>ʾ��u똏�0}��r�\�6;��2.�o��<e�h��#�v܂�dW%B
Zf�tA�>sc��-;j��Zݏ�c���%��G���^��T?�]H�sθi�2�ƃ����Xu�V�j�?9�u�?�x��زms�_K�3��9�rBZ* z��(; ����Xer��hjǹ12*�`8���ճr��=[��	%�����>�!�e���ꦦC���ʦ>���fo}�����˄�0�Di����C�Į��a���WwG4ظ�D�@l�)�C���t�nr�U+�@���L)��K>KY`��iԧK��.Į���J�5��٤&�C� 2I�W���0
�+d��~��j��	�#!�@؁���YNz�a�©����¢7~��KP�JW& ��.�Я����z����\v�'D&�����8;��U��϶C��)��!F�@��3�~B�o��_<Zs�`�j �){$��{�C����Я��oƠ����8,��ꠔ��F��EL��O�����J�+m�0��$�B׎�<4y����9_�����h2��2t�c��86�P(�Ei��Q�ؚR+9tr�����|`H�=��y���dC�zuǞS���m~��S��O8�Z%���T ��6m���ιZ4fƌ��Z澀{^�AG4H��&�E��!�Ջ&��l#���0�������|�u�SЌnEk�Q�*��+�m%�'�B%k`3<Q^B(�����O�c�C���/&�Y�?~�s�cO�m�~*J������\���8q��w+��]{��?Q���,G�t]p�,�dҬ��������L��7�c`���N/3�A�	���1�`��B�7��,w���>-V1-�o0l�E�-�*�:7><-Y?G���FT(�C2�}k@�#T��R�tᐜ`�A��$[w���鉌7�6�b'K��8y���[��	Q.;3�8����ǥ6��	����d�릞�1FN�
� w�����@q��̌ڋ�x<R8�"�Η�1 XX�0���	V�D]q�1QɚGjp���l�A�$��)�I
�B�������id�++��lƮz�.3�J�|W?�/�T1��,�o�20r��u<2U��x�rl1)�~q� �9 �uykr&���D�Q�������7Ε�昚
E-��-X�g?��_�3�̩����7L���nޡ���a�xgd��M�ڧP��_ۚ���BW�BF��H��U��a��Fe�R��;��̏��l;Ybv�4�)�7?��^t�#�Q=�5�ȶ%���J�ۈqk x��ڮ�heEyH���R��s�^�!�x��R~6ه��F�®ц�f�ܱ I�� 7Q<�H�VQ���$���W�=!Hץ�D��:����� �E�Ոu&[R>hƪQ���0�~f{�XT���(jѮG(�`y��`b�hI읥�!1���|i��#�m��W�~�S4��\D;:�镶Lą�������Ȫ3�0�$P+0a�fA�{�a����rP�.�h�(=�{փ����x+���F�I]���u�������S��:j��� ~<_PW���ac�X�롾�x����Z�ݒ��G��!����Oq��J�s�C���a}z��p>���w���'o)���s��@Z\�M��(�ypl��b�U����b'v$�7��z�	%�;z��WQ�G����q7�&a�:��ר��^o&Kե�����bC�b*Fa%�P7�%���X�:l.�{TU�U��jhqCВ�IL���R'�{�g���˘D�v�@+�:AIi�G�@Y ��J~O�g�-��z�!=\@
C 4���u�{RJ��c�|�y=H9S�;�pW�������˚��(��ܙ���� +^M��B��t���l�]�̴�9.��#偦�����Й��h�L�M��w�^��x�.��f��V��
i"];u���f-�_A�c�~�hP�~��ݸ�:�Z1L�\D��9?4�K���г1Ϙ�K�?YsR��)&�C�����Z��L'�NL����ڟ>V�(��	���R7"���MDɈ����4^p0��So���p��4�Y��޵Y#<i7�&kF�qu��\�O�?{C�p��cMq���ٛ%�qK:4%�ݩ�7���Y��@`9�3��}�c2**�&$��̎B�zH����^/GC9Y�QX�2r�Zhd<) PWc�ߛ��	��P���D�\;��	�2$�^�m�?Dh"����h,g�,I�c24����"dBMw�F?HQ4�t�4 �<����'[b@i����H^y7�I�t^�:�M��F�Ҷ���)�͞�1����X���r�؏�	�?o�ȻWcJ���4^:�n�D��/���+ܫ]�*�o�ע�gǢ4D��ab�o
���_��*�νȏ�y6�d(���I*�. ֍�N���b���mS��`8q��Ŵ�sU�JY�G��}���Z�_ɶ���N�X���������2�륩#¨�(&]#��	��G��?�a
`�aT6�g��<y�l�:�{k��y
�O�3&`Bv��Á4���!0�ebWL�+s���	���"�VYSŧ����DM"�|(ו2+yGe��t�0��/�Q��V��i}b��`���i��q:�O���<�b�B��ګ�=*��6@��S�!s��������<GX�󱶂�]���]x c�P�Q��ܞ,1����3�s����4z����#wHk	�//Xc�T��tpRs�+��׉��
��=��듡���=��)�:1�����������4��i��0Lh~�i��1�\<�Od�85�311�G9���H��~I�iY�d:��o�Fazl�5fA�gc���d��v��jHYa��^I!�_t�pnI�Et�-&H(I���7|N�q'����W$M��tȑ �{?�/�D������;m�=�vq	���>>��^,��Z|Z�����'�b�e�60W�o�:V��B#���?���3d��slfͬ��/�Ӌ���*�;}�OK ���"�������ҋ�:yH�jO���Jv�@��7�F2�n���,mb:�h-Y1 �q/"���S���~�p�-�0�Y�}`%���%@V����<2-/؍�ϙ�h��c `=�S�Bl���"��g sVTbH���$��?�铃���:X�F����jX�NW�D�>�=w�)P;���3O�F���r�1��܋�"�Ѻar�����6�������ˊm�n�5�Sc�]B�yS&�� Ξ g�����l-���������:JuE����L��ܼ��4Y���:��>?%�dRFQ�)]m�z0�Cϼ�W�4ʶ~P�o�]�౤Y$��f\(��i�x�g�'���`=Fl>H���w�Th#ц'N\�^�@Ɂ�
7W*��T��?a����?|��?}�S���hȟ%_�֭��(r��,�4A./��W�TzI8��?f�s�I+��M/X7�
���G�Y-��\0r��T ir�}A�f�ƾ*YE:K�הjCH�}�j��禍��`�U% ����;eo5�e�6u�	3"Q;4��9�<X����z�#�iQ����k��*"��D
�d)�Y��Uj���Vo��8X$�LV������O�m��~Lnd�u��
��D�����7}	�5E��{�-����9U-] �H(�A�-PF�1�ߠ��qk�C��	e��,Mmδ�v�E��d�vy����g�d���ΈBITj��������μ+��t�i��r���`<�� ��Y%=1���/�X��K��s��F����T�r`�k�84h�K��S �>\h�V��:)�I�ƶz�LI#�Р=��o�L5�b�� 	��_�ڒ�4�}�����Kp/�Z��F��S�}x:3���-9���g}��%<iG`��ق�+�A�-������ّɮ'Ħ"�X�������j�,�m�Q0�	'�F��kw� ������e,���D?�X i��NP�R+�_�}�X��b��WI'y�_b)x#)F���J�M\̓r�˻ٺ�����"9�9Sv$�����J�|����	�S:��͛"@��-p[_�:јX��{�eYt��{�->翫`Sc@'X���O2T�/Y�����(����g�u��������H��IdM�S���1��0��.%7륏>�NB#V^`��E~�[�M9g����n��p��������8�7!��k���Z9�XP"v��߾�Q0��Di���;N�ge�?dH.T�8Nd����T#�JL�ݪ����i�\%Z��7�r�ͯr�6�e��J�n��2t��EǸ�����{,���_�}�G|�g����p>���2��]�������	��h�^��������2��i5��[g�#��!�	0��0ά),m;U��N?8�@�2�
�����L��ա=�"�����ӎ>�MW�:�r��'��cC�r�f��<�]<X�ā��
p� Fw��yo�#�R(��/=F�	�b�}x⯣bg��E�4����'�z�����QC3�KňU�"ݹ�]�?�{�T��k�oE�}wX�룼���J0DA�t�]=L����*'D���՗�Ec��Ƈ l�8��A{�~hm�쿮�璫���]k��K���@~�ܧ��Jj+R17��.��U?�v�y���p8l�v�BJ!�����O�M�k9<UO�KZ���ۜ��k����+��<1��G�z��K���c��8����>%ɚŎUF��z�fǤ%�4�(��f���{�L�ɧ���:�����
���o�+��w��
��o� '�������D�loWtp�9^ʴS����ϋ���>E�w�YǑ�Ʒ<����y��������L}�n�{u����]�g�,���*�qm<� ��qP�y�$�-�>��4b�_�2��ׄm$��F�"���>��l��#��In��3�KD�|L�抦$C��w�����O�(�sq�F�)kzL��43[����q(� �z����d�r蚡=3Dyy��X�!�O$<4���蹶���b�Ws��k�N ��g��f�1�3���v��	0�Ǵ>�S2�^�:��r���hĒ�e�䂑�C��W��y�3^�8^�2��̈��D�r�v^DJ>���mb>e���G�8��~�9�\�P�P�c�9�$9P>J�^?~Jl����!��o��w�C1�ʢy|yš����S�$������v�5Ё��0�[����������\�0_Px���r���3$���u�0��`�~��-��$�WԀ���{�n];�Yg+²�I{%���|�('c�������S��%�f�7��a�zEQh�C�O�O��򕝚������ބoO�勅w������!/8�8$|Dw@�%���!�,���9�m���쩊�&٪��S,w/�2;/i)Jj(�V�gW�q�&4��T�KT���b�ie��H�^�W��۪&������u؞�I5>��O	�����+5����zx�˱�R\��!��b�<�Xs6���4\��2MJ8i��9K����9:m��3�c�⨜�֯,�n�)|�Z7lDr(�d���3����8\ ��B�ƥ�_�@F����"�38��&>6Х����ɸɛsX��zl��\bp�k��0���@�=���6�E�E��1�SD5�?�6�:��7�����=�r_���[������9)��O�EUn�\���J�/�����<��d� &b\�w���r�I�+A7�l��$R7*���+%�C���&�B�Z;�ֿP��!����Gf��n��M ���:�˟�Ͷ��-M4'9ĒO�&k�:�Y�WP�,	aJ攙��+F����ܞ,Tݘ:�Yt/-Q;���/P�׽�||� ��]	�\Q�Z��6�w���jH_V}y#�
u��p�*Y~���l�&����_��,����2�%@�L�oh���ǟ��;�么H��Y�ٍɒ 	�Acq�	�0.�U3ɹ�TQ�	��vȺ%�Ĉ������$����E���2"���<4����|JG=e��B^�$raltǏ]�Rp�[���K�I���v�`t\�鲷� 2c�6`ɨR[d�#ܱ�r��&r��=��N�W/|��qfIv�_T�ä&ߧ�+47Ȳ�=����/t9��ٱ"�J�&�`Z`�w��3�k�U�mQ����3'�gH�k%��R�-0�F��gA��������;t���h�1E�Q5nEQ^�9�gLHgp8LHX�#l���'����w��:^c�[mu=��������I��#Ўk2q�4�{�v�w��h0GҝW�t_�o�f�-g�3,�'��T_��R42��h�N�]|�����ݏ�v��F�d!�ǭ��o���93���J��N:]/�>6�=f�ퟖ�փ�o4�u[A;bwH��e���V̧R(����v��t8�@���&��_��,��-d���u���ݛ��`5�"�j������g|D�$��<��PE�G)ZN��:Ϊ`_XT����z�ؑ���Ȟp��n�o �hI��+�UI�}
W'EZ´y�E���G&�h�Tf%���yG���3�}�t_vq�Zҭ14��Ͷ2�K���
�(%��%�O���:Yl�X'
�`*�ٱKbG>�%���*�T��5i�kBy�����CY����:]&պeyF���W�����I�&"�^ڳ��ѱ��E0]e�7i��������7���Xu)2�C����T���}C�	��pK`����� �	g$���a5�G����>&�n��O"�z�\ތn��L/o�*�\���c����5_V�� `N/|��m�U��"٩%ZG�M���G�'�=q�8����W԰gE�N"��v�t�ǸW�Rw�7j���}F��m��d.�f���M�ë��,P�7�h���:����OK��0<FW�A��SV����ֲ� Hiy��}3��v�m��V!0�K5{`j��b�脓�I�3S�:��p�8�7�R����b�~,�N�W�_���B��'L����
&7�^bIw'N�����Uտ TiSs�<W��
i ��{o���4���DB�g�e�t3�Â:�"yx�c�{>������7�T�U��1��/~�yu��Ӻ ��&�0!��<N���Z
Y5l8�m6���JS�5��t�J�ߥXY�m� �x/ൿq��l��G�5�p䜓�
.���V��:`���nJ�[���h�����t }�j�$�N���۸	�� �R�TN��q_�����x��B*�'��
`��5������T;�����V�H�i���f�mF���28\=�R��q�Ŕ��EI�,L��P�b<�LS�KE�55�k>����>aC���$&a�P��F9pJ��'Ჯ���s�?�ZF��:3��D��:P�31�����y��iD<�وLͺ�*��Y��B%�H'A��}��@�p��^q�������l�~�Ϳ2SU�V]�]������%1އ�D^�*�b�U>��~Y�!9��b[��!������3L��e@ť���!���%t����)]��� 7�1@�F�Pݘr��q���q�|�1t�jtN�M|���ۥ�D.6�4C���XN�^?����*����?��L|�j���_�L��'n��SA����PYs�b��	siſ�h��OO4Mu�~�"oT�u`������$B ڶ�x���$]e�,�,T�X/p��iu9wŜp� ���VWs�����>�J��u�a�}����Fc�$�Ҙ��
��^Jx�3�C��d-�MX�+eC/��Ji�O�2��[����׈���X�NY<���s��Փ!��n�̨r+vڌ�"���ΏY��{sD������o{�w������9�����l���c����K��K)a��|��s��w���B�*���ؕ�SRE�F�wH�U�[��k�\5�p�߆3��S��[�n#ZT�]Ohue�4��uؘْ˦���(H]�n�_�x@�/���D�j�D����G�i]|s�A<�t��i2��-y�?��R�۸MGf��Kn^~!n���V6HB���n���M5���%�-��^��X�����j"��drԅ��x��� �11'�uɄ]4`�م�V.���z�ٻ�(��a!1ղLz6-���X!C�s�<E�*C��9g��˹z.ƾ$�n��}�)��A�0��F(�؛�x.�K@�Y��	lO˱{�E�7O	�
z�H�ܔ�"�ƕ���*6�\��|h�qv?8b�hbG[��w	�:ͤ��`����7T:�ǣH��ԏ�+ �D{���
^���0q"�c��06�on!��zG ��G���m;g��j�e���JMj��F�d���T܄+��,bs����4��bd��D��w�̨YB�Ie�KV�"�)�%-���� ������5]AW(�QgrH<��J�3�t��ס�:uq���w}�|ף] �$��3;;��o56�#v�rK��|�W!��\�ԓ�#c;Օ9�v�r��T��B�c�]��۰iwd�!a0��-�Y��
N�Pu���c�L�,��Z8�T��G��a��D,c��Z�S(����B�
��(d�Jl��>�缶������G�J�gz�X���ǍݥN7�s�m�@�j�-�m���$P��5�K�$	�5<h���H6qUM�u|�1���J����SG��F�V������=jc�Z�#�d��!�w-D>�>�J!:Dx��(�����gk4�����l��Z�.88�C2D�����knZz�B��j�D�0d����O3����
��+���G�!:CMv��|�D�H,�������oR������g�f����O0Q�L����t6�{e��|�?�.���*���1K!S,)A
�wny��CcB7�ף�*
5�2�?V�	_;���pr�C�j�	<{^��ͅNL��Dx8��.�9�4���~�9���g�~)��j��SZ�G���m�� � '^�~���X�q���۟�$g+Ɲ�T�F0��� �!��+�[R��f�m
�<,�c��I*�
}��4B�� .~�����8	�\�}6�	����i1] ����L`H[��J�t�#X�
�蹾�7z:���y��+�l?Cڏ��.�]��� S(��z��:��@����22d }�=d����ΰ�6��D�t�J�Ќ8�B�S���=
;l�32��9N0�����i��z��}CʖP{�1��_`���P�Zu%��~��+nu ��[�E �;̡�.Q��g��Ӳ8�*��%'7��F�<�.WkX>ֺ�s�0��5%oo
eП,�P��G5��c,�/�6�j��^�5`��'���VQ��s��$�x0�4�ݮ�*�8\HtT�D�P\�gkw�9Q��)Jo��W!�����$�;[�c�֏���敔�j��X���G�Ru����`�1�0ڙ�Q3���q���*���E]p)bm��ۛ�8� ����SH��G���E_��L��<�*�vs){�,�/�*j�@��5u�#t�d+�D�!� +|��q>�R��S
�i+�3D�o����Ӭ�w��_!����I^uo�:�ۄ����]�/���������yd� >heq3����я:���\#�a�Q�#H�韨��G��M+޷����[���(�f�X���je��	6y���#��	؟@Tp�`�J����ľwF��7�>�K�*�yx���BbT�[���eD���s�jw>Ir���׼f-�f[ 
uˠ�''O�"�O�!?��qtm N� }-t-��b�T�O�=1���ws�n�hs�og�\#��CpX��*���y�"i�r��T��@v�FxA~��a��%��D�ES	�đ�R�H[�=ˀ���Ք	�t$%�4�ꚟ ���9*���J��Gq��Q̂x����8ں���=W0^�~�q|hM+'7�P/$0f���d���;TR�4Ii�7���b8�!�M+2
E1�r�W:3�bPz̏�3�VaO�u�
^��6wtč4�7֌p����,ʶ�e�o>���*�9.cY**Ӣ^�V@�>7��a�k��:�Z}��pi�!R�Ӡ�n��E�Ǩ�b�#��F��B.Ϣ)b�\��ܜ�g�5ޥ���}�-�Ao�j!��d�D�5�̎L@Җ�ߒ9	yx���I��`'�k�G�:I�ə%7Y���M�DޱyE��l��"La�bό���Ϥ# ���<q��\t�!5�Ϫ5��Kr����E��w{V��>�i4%� ܭнM�|�_��6ɓ�w�D�_Ƭ�k~EbA�^�9ҏ�{��U(���oOl*ń=���iQ��'%b�N�(]9��2���y\a��f&��\�itz6��te2c�&��Au��Q��޶0{�!�&���ajp�RC+Q� ��h���E>�F#��\(Ԍ5���LKn�Ā'J��sg/�� N�4~�!����8p�p˾X���W�E�X|�_qQ�PٸM��j�:�U����\x� �ýk�� r��ŀ�j�>=�7�hnj�/S�0�$�;=u���C����O�-�륎)VT�[���ܱ�T(���w��014��؃��o �j�A�X�4��I�OA2��܇�ԥ�=�u��#)fM�]rL�5]-`px�zw��ރ�2fx�!��D���I%�?ٞ ��+v�jK���7�I�t1������(;���b��E�p���j���8�P~f�{$�#�U��I��ks<I�F��@������|T�ݾ������GG� o��-�<�9�A��JQ�W2e�`���U���fU�OhXB?����T8ũ�)��Oza�f�|zp�����A����;�o4�(m&*��t���r��N��7�����^��_�#�$��hލ6lύ�J.��f�hrg�����\��};W=�֥ސ�x�_ЧL`V,�1~a�_�wt7=����Zǖ5�a��
�F:�M�텘 ��黍�a�Y5���VU��nF�3��e���r�_���v������0Wn�χ�y��=� X��NV���yH�4�Y�!����Zd��ǯ�}x����k2"����:V�,ǃ���T����<BSL��8��"��j�6����x5i%^":�/��
d��#�9u����nEd��1�0c�����*\�և>�~-$B�:����9���Pі���>��<^��N�; �Z��c�\��}�eY�#�[c.��M}��l���I�D�����x�
�YrS5�M�P�=	��I��f��C�Ŷ�&�RU������>%Ƽ��W]S�ܡ3PE-\��p�����+XJ�ݛ�`��.>��72U���`���X�ެ[�/��P��an6�^���b�����:U������/�Q��D�q���������P\��S��������8��}���4�'P�wa�I�	�1sh���������\X*��5*��'.T�ZvJ�[}��������l/���_���t1��k�zF�F&ڷ
N�g��.@�Y5�+�5I�kNB���CZ�AglZ����[���*W�]��:���8rxX�7��Zfg�n�&r�4.E����Pu�'��gr�-Zs;Ms�č"n"O�ʑ$m�v��O�tQ����2��3����Um�H�-(ˆ�ܪ�MS��¹7	"f��g�\󆟁{fm2������|���xǁ	A���=B��9�k�������R�g.���u ��0�]]l>���o�[����<x�4�0����%s��O��E��鳌1R����U=������P�D�ƭ^�2$ea6�X�g����O;��wDac��p�Q�_q��^m��]fN �J+	�}�n!f���d�ŷP�D��ՙ�n�d0@䖇)㱣{#3$���x�K�)����o��n&���S�"7��=���ܣU����T)��o�[T�(�ʟ��g*w�Ю�"��e����5bh�
k`#ܩIGAd	V�K."����F`IgWrKO�̦�Y�e4�j�	/�T�#Z�*�ѻ����lNq��c��wk(��Z��Ww��_.�^|�T?
Ȩ���U�)���F��'����v汃s��TB�h'�<�ȱ��a Ep0����o�*:�����׈�z�,�$EIŌk�0�6\8\�C�>�7/����|g�&>�0�S�Q�����Q�1�2l��p���%`�Q�!p91fhu-~\�����`���L�N ��_�@�?y��*���x�و�TƖ��Q9��`\��VĮ�ԕ�K�����0a���9*�g�(�*h�Ob��q�[ �*���Op��p���['&��C[,p^ &�IվdR4g1�~|�~��P}Ij6�W����̚=�9�4��$�����;'���w�KX�-��@���d���O<8�B�{mw��y�Ɯ�4׏.��`��"��Ȍ�#�g�u�Ý��{a����A��o�=��c�B�$Vb�2��P=�'E�9��j�������¹�_�:�{���a[T�������+NWL_OL&�yI���\j��h1�l�F��[������@{;[�l��%���cw���p)(�PB6v�63!�]�uN!����K�;c�(Q]���r��[p��PS��D����/�p�^#�a�$��H'&�cMJyG��r+�j4E�[<]���Ie�P׃S�8�1�\Ø[i���A^����<��#��ƻt��&��s��/�7��.<n���Rϵ٥����N Yu��l����UFz�x��aG�sd��S5<�p�\N.}��ت�������US�T.dJ�����B6[qLׂ�?�Əv�X*���)&ɴ��}L�x�!�ox~���O�=�HN���v�Y��:z7�^����I���U�P�)Ǐ���{���`뼦�]�jD�e\g�BH���>��Pi(U��Z�a��Ȕ����&�B���������kT��=~R�NQ�d}[ a������w"4�[4�U��C]4���	����|����R�I����pF�z�	�	Y�����U�'EG��I���Qa�<|���!�
"P�8dkC��qlhL��U?�
�ƪ��.T]gD�8��)��2s���Hݦh~��o=V ^]R\��M�Ά��X��F`9f��y��6�3Z��t���d�9�ݶM�i6C�0,'sf�rO����NR����W��Z���ms܍ӭ��*�ƽ��x2��5R�M�_��hD-'�^�V�"�[],P�xrBV��
����P:���X���Ԇ���c	�(ZΚ1��k6_��.5�^�O^Sh�J�L̋��s�^3�2n����3KN�>|u|i�>	*w?����`_P�e�[C<�
/��/gz@��>�Q���p�`~|��HŃ�Y�qj"�P���_-Dxo�������!��s���t�m��I��7��K¥ȣ�f���cPv[z�h�ǸG\��V>�Y�k�K�s;U�mW��!L+���e�P�&��g%�H`�!��rN_+a�p���˲��"ߋxx��]�h���n=H6u��F.v7��R���CZ����?5�F�0�h�!��5�(���WBũލ�j�iS�<�đ������� ��s���,�(�J�,O%������LE'��3[Yl��/kS �f��X!�jK��jW7KȂ�Y#-xAQ���fL=^b}[^��~�$Fk$%���9PK��#��&GV��Ӵ��
Q!���xP��TA�7&�Y ��� 
BHs�TPU��}f���?ы2��j��*tH	�[O9h��X��߃��{����zt2��+�AJ�(HV�C�8B�S�x)J<(k�����w�J�{il�֛�����H��nTK�B���$ڧ �Y��D�eO�P(��l=�-]�}�CaTK�O�`�X��s��'�SJ���7|���<_^�S��)�C�fP�ũ�8|�2r��[|v����h_�`�6T�
C0���޸���Is����dW��Ҧ�/�#̡�O������$�ba�4ʉ���=����V�-3��3�s
(�CZ'a��Y0���3��a��6�,�C�B�8�AV�8O#��73A����5aG#�gxYE	I��0�/̅�g���9O��II�F�PSE<\!Gy�[ʴ�E�����1�O�Q��������U�z�a̪����UI.{�s����MGs�дO������\P1�`�@T��v	�E��hOg�p�?�'�`B�!�v��2�}�ZJ���i���~�m�av�M��'�}��I�[9qA��"�C���muH,��<������er�'�*y��]��b%q���D�I�h?+�/\ӀU�8�YP1��Y����qq���|��( {���=]�q�w�-G�i����u铖���EE��};�?l����k1�=@i�H��(���B[�v���C����h��$3ʽv ڪ�WK�̈́�,e;�Gb�OH��[�Y��#��w�n>1�v��=�pg��=_ə�<#�}G�c#CI��ӛ�X.�5��?�d��K��[������R�%���V,��?��рp`�Ίt�����'�G�"Pʥ�s�g���M�;?��\�.�ͳ>�s!u�!�V��m�j.����dr��� :�&En����9�)��[�_B,��qL��N���
��0Q!�����Zq�ϙJ6S�+aQ-D��0^I�x�0F�p�&��5֙���٢�ѽ�B���
�A ��O��v�1
5���V�2�j�r�f�* x���l=t$�|�?p���\+ޤI׭Q����,z�S�x]�b��b��q�h�lVXRGtY�D]Ow�8�c(af�ӕ	�\[�M�c�6�LR}ZA�z�*2�
�?���$�EK1�g|�3��o��ߝ!��V�j�5�#ܧ�,z��rT��N�e�'�T7<m
�Lֿvͩ�6������2��2�0���By�}KQZ;�+����nh
2�I��з�H�6��CG&��ƛ"����k�֎�|L0�]�c� \���I�Jew��p�����{Q㝙( ���.5\_t�c�^v�` h^��I��lg���h��'i��3���+�Y��y�HPO���3K��p�':';��k�	��I@�����$�o:����2��w<3	��O�'xhXz�0S��-�O�כRK��<s}_��ؠ�G��l�,B��98���`�P�"�wtV�㰡����\��`lI������i�Ʉ����I��#�o!-�ī;��Bs"ǂ+x����7���$���P �J����}�M��eX�.M�~*�z}Ώ�ؖ����o!M�nx�߾h+.�D䱉��g�@%<)ɐ�����r)�)�\J�\���#
��q�*�^�?�ߞ@�M� �������[�~ύk)�#v��)2u)Ѹ��w����.����H�br�$�h��V*��F?p��CC�q_S�j���n��)�3�HM�?��w��\%�wR���xџ���`��P��1��b0\j]6����n���<���\k��Wd���$��m�n��6
�������ʯ�����&:���~M��S�{Y��eg3��B��n����q�Cxv@��
NCǇpw�'jƇa�,Z����x2���
`<���r��,�S7���U�1�{u�b�UQXp�k�#z�N{���09�&�!Er���v_�;>_j�GlD~��U�%��=1k���G
d�NNl/��EI�/��F�x����������P�JY�˫��p�!a'�o���k�)���i�e��^�	�蟵���[�n�]JTζ)�z�8�4A`�\[���dK0�D�<"��<����iF������n��2e�c�3O�4����3�~���xb[W�<�^f3�P�`ǁ�Q^�j�$���8�x��_��	U��p�H�����6L��L�i�����5�c�c�5��ޜ�U���P��&:�����a�����Ⱥ�x��'K]�K�GR��� ��(��M��3���2�o��s<m��V�'�b*iW��ӡA����W�Q@J�8������OΛ8H��DX�Y����U
�l��=�H�8}{���6p�l-t�K9�օ�!�Ȝf�G<c�!�6�0|�F�7�T���4*5���F�����Z�����ȟH�Iuʤ�0o �_����c�����]��.���<W�e���g�U~�l滜�?Y�=���l����+�yw�Lzj>Ed�W�]�&�w��0�7�U��Q�YC̩e���Y�Mn�`������r��A1)���^8aG�L�C�cT]qW��
�w���Q+jd!c+��zCF c��8Gݧ�H:��Vd�;���@NH8���g8�_�}'�)Ei�s���H�|�*��	)�d2�i�0%R��u�s��)�a!�R�ĦR� 0dFF/�rk��O�����Zz~|��+^���ӛ7��%@���V#?�!�R�^��	�*�8KD�8���S�t%Lmpc�l੄��N�P�y_x�;����i�������-�}��BA��W��_sݽ������3���H|�2�v4'��T 'G���I<�˱ Wb�zb6�!�B�g,�z��~I�i�)�+�epmS7�x6�$�%%,�l�ҟ���>�缝�	=�����{n'��2_B�F�b31}<�yS�z؊G �,Wg��H���f���+Gs9�P�߬�������0���ڼ�*�	}�6��<\K̝��^\-U���i9i���6$"6Du(ļ
�J��>��
Ҕ5���ED}�RȌ|{hTR�&����?>~���b�x�f�A���+	ƱEpx��3���_B��V}qs�̭��p�h������D�5�M9Ir�M�i,~a#����9�o%��B��q��CS���k�m_kS���9s���	����P^��S㢠ƾ&$;�pz7�~���s>>e���Tb�Y�i��^�M���9=�	��CE�S递���Kޱ^��y�}���h���v��Nj�T/��.��I��D�K��:��� ��,��Ntio�����A�|����!ĖՏ�}��]�v���p��aUp�4>�P���[�0'���=[�	�^�G�嘳?%z��)�2`�d�C�b���U/`���/l�����B��2�O�-�t$��X �)��@�@�D��@�@�rܥ H�s�EZ4QJ��m鑀X����v�4���ROF�9O9�2����/��^Ƃ��@Mv׆g�U��7v�fՈ��d�q@�lNq�(]Ż�TR1����E�S}��mE봆D;r�n3���S��CH]��Pվ��Yzx*����ʹ	֤�D����;i���&Z�O9�Q�JWQ�`V���mA�m
[��.�5�<�����l�����[F#���̨����|���?U�K�?��5wQ���Ɇ��,���!Gմ���X2zXm)�$L�cӼ���e�Z,)"�&�g� �fbU2�ƅ� ;a���j=î�N-�='�j���~�2�>/�'�ρ0��F7�ֿi;�州�+�w�nje�oT���Ê�2GJŘ�`#����A0N!�Ug,6����k!vX<}$c�ܢ^�J�_
��;�
� ��^��4%���� ㏶,���.�iD��;s���4�k��9ǚ�7������C]p����_�TlhRL3�խ6Lh�G| �_�$�Br��S�׋p�F3��*)'�zʠ���2A����Bb��I����I,��nk�	�q�����B�h蠑I3��+Ѭ���o�B���]F���SC��"H@pbI��b㟲"֙|��#HǗ�<I/u�%�_JF'	ж����a��_�U!�� ��?����$��V���8� ������,z빽�[C-��s�Ƽd�/�����/�6�l����Z+0ɶ6٢��ӽ�yG��B>�A����UýT��p�M�7��ǉ?�����0��.O�vo�t��j�z�BR�7re�m�N��{#iTH��s�
���L�E�:g�L�+z_�[�O�kUQ�s����8����̢C純.7���OK��������۳
ǎ�e��Ix��/��hۛ�G@��H$� ��F�?R*�e�E)���1'y��G(�&�%	p�]P7ez(l mh�Sw |�
OdHCb��*+���-Y<�P��6t��TQ��)�=n|��R�)�~����}K�Fx�Zh�QǷQ����P~K��F�j�b a��Km�=�bJ �ؔq��_Ƕd�N�����G��?��#�^V��X׺�禚����Rϖ�E�C�IM���"uh�=�9��T*m1{3�i,�k��-�GB���[^X^�2��м���Z���U�֚��ª*�c��Wd��[�E�e�d� ���K��%n;���ȣh�^�=�
Q�9��ؗ�:?�� ?c���R�v�N��"]�6���C����t�BOQ�`����Б�����,�e���/�[���1@����N��[9!��N���oZ���.�>�y�Tk�����o�dU��օ|ؘ����&n��zGN^0�Oz�*B����v��&7���xgYwQ0�9�a�CR\nc�f%���'�F��Bt�������!���X�����p�Hǜ	���1$p7�o��9���en��Q�M/�й�鿋˿��^c��!ZQ	Q�>xr�@ѓ89(�Iۊ%6{z㲆�c!/J�f*�as�H� 9�<��\Em�����~M��#mH��E��jV���K��.��F��[J����C��?�|c׆9=��~�(c��q�ߖ��&<K��u��oh�xF>�`gǐx6�7Lp�l���W�G�#$�yҾ��JK&�N�[#Y��-���P~V_��P��-Ar��� ��F�>�4�7�?����"�r�2�$^��y�+�Q���~�����.�?<�3оⴽj�.�,�D��Q��� ��"Sq���J�ޕ��y�p7zp8�:ØV�?��y��;.D���Y��KRg�!Q$������gM�������~� �Z׸.�b�ԶBLJ��o��K�Yx����~���B��7g溵����i�lVm�CS�v��݁�T�� �k�8-�ԇ�z|V&cd���5���9z�M҃����]���>�G+�����+�EM�[�`.2�ؼ�۪[H�V��6�*��>�u��4��v{�����
���E?H��K�[F�QO�~����Ĥ�Ču�0��?yc>T�E4�LZ�߹��$J���(���yh����e0aq��B�z����W�����φ(�l�r��Ne�D�Kq�vF���@�xq�J�D.�E5�n+���\�>�n�/(��S�z?�F��ڤ�%
�t�{�0rE���-���$����S���A��oS+�p�����8Ӿ{4�#�����	t�!�E�t<^E�ς�����,��~r��U,�K>%�@��6��@m�@]P#�\��H϶(��u�	d��!�k���0?!ZV��@_�
"U7L��!�ؤ�e��W^�)�]&�:dČ����@#�k#�e-�*�iͰ�;l�#�풸�p�!�S��L���������9� wɊ�MX��]��69��
�-����gX���cu��B^��cH���ͽ�"p^�;��Jc���Xǩpᫎ8+�h�����e!"��ri��dFG�#�KYI$�� :%���xU�w [n;�-ө���. G��lli����_/�>U|���w��:�~��D�-�<1��:��c`���3��,j4��a�L�fw>U)�%�?]<Tչȴ�.4��*K}�;�M*��0�����s���Q�sQ��FR)V���� �����XNeW��N-E���S ��/�=x�*�} �񺝍(�ث�xd^F�vm?:Y�g\�H-��YBL}�vDMM���8��vqrrpߓܶ��"KV>�fi艶)��;�;�!f|�Ʒn[H �)�ց�o������ޱ�:@t��r��%�=4�RI���Ґ�%s���أB�ѯ�q��tz�y�
�2ʅ�2��ڰ�+w��o����=֗���M�u|��y4�[:��c
f�0Cل��� .���͍��2!�tU�Ђ4f����H7wz����%�/D���$��J8M���;u�,��.�����q{�-��H�U\�)X��[�E�5r��RM(&���]S��Vf���c�9�'� 2lpP'�Ԥ���ܖaU.p���2�=����4�E*2���j5����oX���z-�TY:xK�{�'�l��yn��>��li��y0h���0	�����)��V�	��,��P�ޞd,��I �@b%l����6�Ht�,x9�$	*A�.N��ţ'h����1zyA�C, N�e����7_�ucV:�}6��L�I23��x~���d����oY����g\�E��Ca%��4@�֨�E���ʨ�?+��Ñ��ڱ�gWV�Oڬ����W�-���g�>�hܬ�)��<�<�(����Mi��ggw�5���pȚWA��,-L]ȫ]�F���s)ϼ_��?ޥ(ƀ~�oE~b�Gn��������������lBP�"<z�(o>���1$�r�@�@��L�:���w+��0O�I�
��U	;�a�׋� ��-��4SuH��"�r�*�0��o��[g���� ����n�d�������#��_Ǉ��/w�[�B��J*�Q��m!�`�tH;�U��V�,؟<c{:�O}��DY�|�&X
ҒB�ۃ��"��	&*��_^�	GZ�R��_��P�w�����	ax��vW�ъG���ޫ}��P��g�%�a_���)�l@wP�7S�+�eA�{�'M0�M�)O�{h�
�D�yLS;���6R�S-�D\H�O���5 �@�7��<��\Lq&�re(�q�B%����"�[ad�����R,�V{���[i�;�'���Aq�f�����J(����Jm�x�����W��&�5ř�k:ӺN?2~4��$�Q��H.&Y_�(B��@��8`%a��fV;�ן�U�Jmg����i(\�J)���dwo�
���ҎX�7��^%=���c��WGd��0��=�Ec���Go��?��q��!���vdm�v�&�u_՗�ٛ}֮-!���x�`/���s���/=f{�<;��1�q��~c� �Z�8�)�, ��-���}�4ݡ�L�f��d��K* j�G�%��נ�E5p��S�߯���Ɏ⚐n��%m�ڞS��6P�#�w���������N����f`o?*�rRc�м3r@(1;���;1�P���|��H̚����P(eZ|���MNԼ�U���΋��G��#Y4�2��I^���r�mSH*\Z���jx��S �dNڏ����jU�d��ls>E��b����L��͸���u�7�K'�%F��}%h�(|6��G�q-���ţP�m�m�%�����{S�*.�Ǟȩ5��38�~��I*z}r2�_8��Ha7��Nw�'�9}x6��8���-ј5�M3Y��	�`u�n7gC�:J��MǪ��wϣ���=n�ҏ�A�n�W� �����D��R�����г4�e�`��;+�R���f�U�h�3�6��y���'�k�G�u
�� 
6�H�E_�~�4r�^���vB�n���E�)��V^�[����/�	��2��Cш����i���	�M��-��n�ґɋ���_].�p�Z�������p�����C�Ԁ%K�I��`&a��em�� #6�b���x80UR*��n�}Ɇ��!�l'�&�;O(��ȯ���rZ�i~�|j�Z$��k�R�tV��Z�.�3��F�2�i�����Ī+X0JY�G�@�� �j��M�Ll��Gx������X���TV�.�q�eʈ����0�a��6hbc�4��+F��(�^+r��n@��3~��?�tSL�_�,�7\�V��2~��'�3u�Ê���L��X��[E�ĝ/c&p�{��
[hrTW���l��k%D86J�}:A��E�G�\�[@{^���ا���u����3]��)^���\�Jwx���7V�
@,((�-�;e��i�_��&(3f��UK�V��mC�x&�A�ڌR�c����?�/~��阳Z�����3���wj��*�^Sf�O޸���Dhv�7�@�t�Y!Q�<Q��)���Qf|�N�W��������j/e����i���9�"��7�u-U ����Yg����Җ���zH�Ks��X���O��"}Z�D�Q\�Ɲ|�t���8��ɻR���CC
�^�G.�p}� x��(���� ��Thx�P�����K@���|@��+u�n���#���E$x�Q!p�x��g����y.��Dy���)���cd,��q�)�:SO�;��2ǆ�=����ZK"�B��a����q����kܦ�T�����u�k|!).1KȊ��T~� ���T|���JhN2ۛ��(�bJ�м$�E�P������F��;�	�D��m���R�L��HW
B$�v���SQ	�=��Ŗ�#��������w� ��͆��G>1DЬDcT�8m�{�I�ӌB�"]lg��i�7������p*K��IXF�HY��ior!7�lt��u��۞͏I���|�F��$��*��A�G��p��3�SV��m8�b��H���:���4��pU	��[|z��$+��1����똩n/X2
hȺ��X�aIo�X��vov:���8;C-fy�ƨg�����Q��I��8&Y3�0ۖ�ɹ[!�2��o�'���SƘPK�[��=>��f;=}�;S�{F�\����UԤb�%%f���`I�TZ�W	�A@T��?I"cC�2�K��T�,
�f����>�i������9�h�Gw�!w�,H��A�.�,�l^Ͽ��w���ԠrH�II��|��/?/��	A1��=%0�Htk�M�sQr�.�$Y~?e�ƙ�1��U��=�1~����)���p܁=5 y��B��q>6Ym8��� l�(�9��i"���A�|�t�5�p�����V���sS��W�������~���q��SZ�3��v��.[
�(�^��lr�� B��i���֤�C��߬+S�RXf4�4�)�t)i��N-���$�Z�`��B}�D����+�4QL�9�S2�%��r�2��pS/8-��c qռ��z�ul=(5���
���-��l�A�w�z\�������٩��YX�N�nB�
Q�kb9on;����s'ğ�&U���}�4uk��w:F�p@�58E���l��M֤6����O�)|2��g��<�ꇯ �!���o|�G�
]M
V��.�Dz��*�`�%�z'���g�>*��}��{�m[�nԼ�̊S]X%��n�x5�|�������%� ��GBoM���tH���	M�#�5����V]uR�s�VA�Vg�O��|�ٹF��ō	Ưs
¨�^�����\"- �H@�b>���#��װ-
+�Ӑ�M�����͐>˓�-�r�M z<ሄ"�޸�a��R~��nۈ2%����U�1bU>�7UԢ�#x���V����V����ĝ���M7YgRR����y����/��Y�Т��q�}k�����C�5�X�t���b��2.��Z��k)�t�;Z$�j�#�w(AY�!�Q�����R)x�51��X�(��m�6��N�*hd���d���"2����f^&Y%��iۙ-����XAOa�����*�i9����!z��p��`
p���ǰ��,f�N��G�.-mŉgGF�qF;0%�Y��%���$�"�F���&��w}��@s�j'�A��?�H_�s�d0L��V�p��QT&��W�n�L_�Հ������Hsܳ�"?�_4ȩ��]��5qܮH�H[���w���d�e٣��\$�H�wjԢe�����W�bGlѷe����a�Q��}���!e���ߘ�*e��u���Hd�x9O��ht"��^w(
.��/*P����(���E���q����}�����B�vC���w���ۺ����K)�g��n�����x��G3s�:0u%K�aT�hr��em�L�ҙ�����Qp"hN���S���Vmx���������E�G��(��+���!0�/P��`9�O���RA��0�n,m0Z:�_>Di�1�lܝ����K��^^�2"�M��ҴZ[]mU1Ъ�Q3}Ī����a"M��q�(K	��R��Y"`%�q<Qo�]�����5�Wh ��p����<�O	����/=�ģ����W>�AsE�V>NE�;��mAR,��$�J��ظ��$6�s*_U��ғ���Y»�ɦɟ�&���/�fn!�ʜTg�,vw����������%n���U���1�������V�d�;��g
/�1W������a�y��7�H�z�DW���{w	4�u�������WKP��j��2��'�~�IZx?�ЃS���}�`�[���?��#��T�D��^ZK��6&���5F��S��=7��@�z�n�xI�z��0V~:e�Uɭ��e9�l�#f��;َ�;�U��{ph���XidTH����+�:����p\o��iE$]�b��ο�z��E�������¢Ia�}�E�.v�!�,����Å�O�Q����,����#t�O��,�A�d"*+w?qQ��[�����R�ut6��7�cx�ȗn�_FOe{/|�Y�����D; ����ϵU�/���a!�q�� Ay��Syj�<��DU���ھ1�!�k:-{���,��@e};�R�u\�kѻ�#s��o�c���/.�ws�O�5>����C)5\�"�X�s(-���F�o�o�yS�n�1����I[��������-�[.�]e�P�݋��7�(����Ɉ/�yϱ��o��ց�춪��,��{�V��%>KV��\���	T��8뇮�ZR��(�[h7�b�2�ٸM��XLn�-�;,:ۢ��^,��V��n7�$C!��ڗ���nmpS��4ډ���X�9Y��;�f^m�&��|d-2�4��ǁ~j��Ӥv[Ӄ_��G��Xܐ��KoD���rC�祼�����[H�����UE�S��:�$q��B�Xx]��P�閥�x2[�:9H�\�B�L�S66�QTi��ƙ�.m���A���&,7�͆^��+���D̡v��1U0���9�l
A��{fg�-H��-���4��a��ᠸ_sy"��S����j��O ��8��=�wt�Lۂޥ��������WeӁ �<GT�p������B�HőW*>UK�P=�A����Qk:�U��d�������v^V��ntUGNR7i�V��gn
9�<��Mz�a{�^:�nP�jlC�vۨ�`�K�u�̓�>eWn���
h��bP�+N��!���D�d�C���P���z0����ҫ� �G�0���ֻ=ӕ�yP�o��^�0�[^��O{�"V�Z�q4]G�/���.��5�S	����4��^p\�j%���{����}�x�"UBe�\�`�Q�-�"�RY�	���;�r�	:�c�s�Ğ���jK�4%(��9����H��9C��-��sWR� w�.�%�?ߏR�����/^[���h��>���m�o���C�_Ӓ�+�e�d�N"^Tf��^%���[���D��A��3م�TQU�g��#gt��\ㅶX vP�[�B`��>F��r3	ܮמ�ã:`a��>����XŢ��~�o���r2g�J��mT�QFp+�0�&a�ȝH3�R���d���j��¿�U���~,`�k'��f��K�Ti��=�O("Mk�"��� �p�؀�^��z����M#-�o����÷��$hjj�2�(ȼ��Q��
x���m�t�	��8���~kt?�f�1���ӥ�����/�YɆ�����IN���6�<�Re�mڊ�a�uί���-�@�O���T�Q�X렙煌{1�͍8�o��]�l�t���%6$����<��E�J��?�0��x�p[��u%���6W�z+u���S��H�燉x�)cj�Sg�!�LxX�߾����!���7��;BQf����R��Jgh��!e��/gh�a��i�̷�z=EY+��t��l판���ל�,adZ�mj���E�r�K8��-V���z!k6(��\����Y�;N��������([��AJ��6�d��^��X�{��<G���0T0�J�:�6�M��TC��v�=�cyy�7
�qq|FzLa]%��a�ƙ��=�ji��P�U0��%'L��C}�?�Ӹ2*��]��Tl4U��S��}'�[yv�g�
����*
a<<$��G-(��cR�_V\<8���'��:�GT��I�i�2u�ؠ�# Tfȅ2�F�]�'� $*-1�ZF��g=�.	(x-H�+X�����6��h�c��X9�k��gM��,^7f�W�Q����=�s�_�Z�*��CN/�P�gcs<kx?�d��c
Hw@��|�� ��Kl���\	Y���yk/뽱_�|���N-(�P����̈_y?�ǭ@���b�c�kЅ���Y��;/��&*��	�!�,�VP#�+z�D�!�m��=:+�.Q�aC�����7�}W��󫔃� r�i�9�+�L&+��������m<�Pe�+�G5j�'yE�M1S��2�!�;��s�Cd�"y6l��4��:�Rg�E�����~j&���w)rh��ߟ�� �9ir��WtU�z2�ȯS7��0fhs��_����5��Y3�GMƼ=̇�}���K�㻖��_�r��ؑ�;��oa�;jƴ���Y�Cg�����r�wѭ��N���S�j|��K����'� &\��/�[��@�y̌X���R�(_�Vg⠗-V+��0�Y���^����׼k�5Е������5����aĊ���$!xb�\�#�U$�OC�n���Lޒ2�6E!긁�>����st�:�Ra�9ʑ7H�l�V<'�z�z��~%nG��pn<�1۶x�殤���8�����=��J�ݮJ��w.>���`"@w^�CyTj�� r����1s���I��#l��8�A:5�![���}z_
��\��9�:�!;�`��z�Y�,�O3���)!�Be7��<w/��sy[�q=��A��ht��,�^?^C�5%;�t�5�����
-5���𫳌���.��������o�_�e%��'�f��_�� ���+���c:զz�KQ�O�D@R�]@~�1y/��[�=��r��`okez�f�0&��a.��l .�5�zh�~4�5ay_P?%�>��� F�߷����S��o�� � �S|�ߑ���)}�izm~(�����60gLMڒ����ַ��7Uc�` Ko^���{8������-�,�Y���z��O�ێ��B��#��A��]���6(�\�5�\�qj�*<������n2ፗ��u7s�zC	|������9��������$���PsM�l�XV�)��@�� 5��X�YY;x�%'�0X�@W^�B�X�o`��7U����_7��j��#��/�7)+�j�_�7���V��M3��<�ŏy-��l9K��45/TN�D@�I�/bAs<3:�t]�Ϭ���};�_=e�hO|��XR��V�c��
#w��F�ZR�B<��9�5OZ�\�jW��Z��*V,5��(3V��/�}�E&]�9D�U\�Q` �(�lcLx�Q����_:��>���]������]���J+�|�͛վ�^�	��%���L��i_Ç������=O$�R�4Q�<"x�j�@l}@��>LoB�-w�h">S�Z����{綃ܳ�A�pLܱ�N���ţ�Pw��?��x��e�*.�?��:a�|sס�V'���2Te%o%���om��CeeX�׮J͌ۉ:��e�/���+p��:>E`4{$vԅA����	^� �hZ�\�`g�p��۵�Z�A�|�Q'���e���C��&��R���,Cv8��ﲕr`'��q�L��O�	s��>�]M�"ʌ{�aR���
\��%���}����o��f��/���6���?R�J>�D��!`A\#?���Ude���u@������6��a<L��b��΂�逸��^�����X�����������KvS�%ѷ�I�q"%(�	�1ԍҏtM���,=�!���E�m*�g�u'`HuIPp���zlh}��)�Ȭ#a�Q��T��8�q/ɴuR���
/��>�x� <[x�
&�3�QM���J��h�}!�V�n��Q���%�n^�Q*\a�o��*��6(���g�e�?gكq������u�A6%�"m6��x�L^���˛\�]�2�?bM�\f@w#7�������מ��۾k�x�� �Wi�2a����>H	�4gk�-y�A�<;�O��{�}r�-U�����nr��]�("�\����Lc��`Na����一��6%uEBSx
5P~�4����%aލIL]"}j~ߧ�Z�p�� #�|ڷ3�(w�VV8X?�U�%�u�C2�97�
�w�(O^d ��>T #�=�׹��B���`k��,R�K����Q)�h�BݰG�;�#O܇�FJh�T�R6/&���w�7W��D��I���t<����ɸ�����%q¡-���w�pJP����ߵ%�\*���'2l;�l���1�ɳ�L���M�L��{���*4-SV��(��C�.��~R0��}��#[������5(-�b�X�Rq]��:"t_$S�|��d�l�^+M�<4��Β�����H1,YJ�KϬ���i��J�T����]�>Τ4��)P+T�*�KXX�L�}Yy*}Pb� E|�}�ٯ�2�V���UZ���8���o�h`B�L���������iB�����f�=�$�w��
�U��b�h=�Q ��o������^���'��>�¼�_S�Fb9�]n�~7�q>�Cy���r��O��8�_��6Ѐ���F�����fӚQ"�aK",\y�a�fE!q�ĆD�ϧ	�������/R�~JI��R�a?C�'����s�����U�V�C0�n!�����z�c�mb�QXA\�B��{�h�zF��հ��F�{�.4x���{f�/P�b�i�?<��ϲ��93�%)�'�TGIc�gDKE؛*�� ��b,5�t�=��-��'�¸ؑ���r�hs�(�uuq�����K�O0F���'��a�����0�@N�f��C,"]�_�D�o�aŁD��ɀ��:*�Y�<��QQX�՛D��-�8kū��H�jQ24�y�Ԕ�S3k'c��W�ݒ��	�
�<��^d������{x,t�<��m��8�'l��Q�;�):#f��S���&CHF;�����3������ݎ�؄0��ۃu1���`�Py���Q�t3(}����B�h��V�o��"5$2���B��90~�!҃o�lnfs�g���6{/N�N�PA�'OA��i��xm�����s���*���/�x�J���M��,u��"�����	bg� *�e���+�����cQ��ő��� ��h�[Gȷ����J�Q�g��
��������j!��$�S�p��3A��`1��3�ceĀ�
c'9����w2��;7cPG�Hf�g�hm[�̼���.���R��q�=��G��&6�h�=�cg���e3ᝒ��I�"6�6t ��_h�ь��yTX������q�u�RyxvO�l�}n$�N�5ŞT����Ȁ\�]���m�R����֝���໥��"Їֆ&}W�����U��sk%�n�cyX�A���A�k�2L�����zxBb��W�Z�EK���z��� V|�']R"�@� J��i	��:�SȰ|��1a	S��:��"M��H�&?l�CTB�GI�S.B3�U�@a��9u�5��g�:�I���^�'[��$b�	UH��M�gX<1��vm	�� _���?���i�l")�c�m� R l����>�q����s�OCF]��A7D�Gȋ.����L�q0- ���f��I#!7РH3R��#Bw�T,���BVe�BQ y�"�m���7s�:$�P�R&K	gE��q�����z�>��崋�6(�K@��S�J~y:�`��M�6��mt�jR)%�%j,k'�M�;��n������
)`8������k��e惊��{��k�Q��P6�̈���B0Wxᒟ�2�R��Q�naEk���>���'�$�۞�[�C`~��|�;�e��8���GXG̓�0N��B[�d��T��Kud n�ӻ�>'��v��q3��g*���S�N�s��aA����7�M����[�UVn]k�����Y�8b �3c]Y��F�����QB���أ��e7�/P!�r�/���'߈�֏�$�_&��{\�bQ� #ɋ ����5�+I.y�	�K�u��N����\X+x�����[:r'ь���{�.��F �IrR�\+8/����R�G���k@��ȏY��d�� bs�]��z��i�U�������ydޞ�K�?������h`��2�Z���[S��[����%�f�y��=����N)�,Ή� D1yI�hTՑqV̹���9^��� ŦS�9�`�S~�Ǣ]R�>�m����7
<���ʡ�\b/��ËH_¹펌�G��i�?�(�}E7/�賚�m��֗J�^�!1ڇ�z�v�'�jD-�0�u�a����h_�8@��7fF�xHfV��,�態5� N���t��Q�uLIz(��0���R��o���H���V����+MѺf�|�?]�(BAj������q�?N�|��б�а����:F��W&*�G�q=)%dL�./t�u/�M����ۆ[�,Z��-KM��r�@�S��N�ݴ�uk����X�Z(��tgJ�?�������ݫ+�(����Ѷ?�����%|��IŰ�o�=��;f%�F�ckj�#H7�˒F_�e�/����k���h"��c�g=����::��J�v���m(=")7}9�:u�!������"�_�4W;װvd�>�#5j-Zi&��Ӭ5!eL#�DIC-BkhG�M��6�1������ˆ�F�m��F�GM^\�_o�р�M����v#T�y��EB!�����a<�}��*+��O��M
:�h���ʧ���}	��iso1����b�$��nw��f�؅����K������ͻ_��jH��;}TȨ2i�۹�9��k����@�F�Z,#7%	���,\uLg5<a�GP�D"}a��c�
�1��H�=�0�`nw'�e�7�T�z��U[J���3��	
z��|�c i]`6 �"1㴆P��&h!��sӯ�@R�9����Q�[�Y4S)���z���9h.�Aْ;�:�Ɠ(OٖZ��߄섊I�F�ls���S�	��W�Gk��p��T��&��/�H�H �� ��+z#rj
?Wd9W)��������`�{�N7�/N78t��������'.OY����rɎ�9q-�,<�>��葬J"�S��Fg8\���LB����!q,�@L��0vXQ��戛��ӛ?T�4���r��Ƴ� :�
f����
NYof��3uh���1Z�	����R��\�T�9�)OV�_C�{��~N�s�OJ.�E��L�� ��׋F�dաj�<��PY�\IX�u��Tϋ�C�I�<�`[6�k�+;YЙ{��}�9�8�	rb�[�E1�G�*�-Qȴ0U�v7��x�}�H�y[�SO����4���7�Z�X�+3�*x7�ڗ�ߤ^�����c�d�~���w��:����`���"�m�evS��	�9���eÔ:��
����R�q!��O���aB�A��{Xǯ��&-Gʹ�so�~����}���Z���txl9�VKQ~�����vW���������+':}���<ȁ���BN��V54�3G5�V(|nF��͢o~�.��C5V�X�?��I���+ּ����Y3���yӽ��~����3����<hӗ'A4�EU>�EY�Ud���ė��Y�9�7o�����t���x�L��/	�O�I���1S������n�a��΢G~�P$f0�w>(*����O
���R�\'6�H�b�p�jp�ŕ�f�B�.TG�%��Ka��'$k�(�a5�N�6��d #������!�r���?�d���5I��*��"W��Sӹɒ�QUZ�T�/�!�?�*A s��qa=���笇��g.i����CNά&
�`��}�/p��Շ�F����A��a儣L�e������@m �|{�򎹘��7(r�k6f��ɷ�*���LHL�?�hw��r�,_A9�ȷߟ#��K��q��n�{QTf4Q����E����[�n���I�^��6�I,�
����e��M��ܨ1fzI�`��Z��a�����8�FK���i-l�������V^eަ�	S��̢(����Z �NKB/��X�/B��f��O0Q!�",��KW���+촞w���%��@�n�}g,��;�t�DJ9!��[��#
�=�P�����9���#����k��~����qa�"�$����b	������V���9�p��ğ�,͠n�H���$��b����?r�l��vS��_�<6X.�"�����F��9\�5�uCn��d��� qC��*;C�MAe�u�Q��n����O.P|�}�.~@'ʲ��<3ʹ����k��|�0�֭�EK�����1���D��xO����=G�d�X]�"��8�7�!���Tl�7�	^�+)KD��z٪�{+��>ΗB�kQ�Uc�U�p����M�ڏd�w7Cd��;�*I]*�}baXC��і!��?��_T��6�&ׅ��,�DisY��yDO����Ī�- >�!DS>嚲m��U=^iz�e,
"�~-�o����w4�+ʳw���F�_���/y7�j߆P�hG��J��#:���޹r���H��Ű���o��͒��|�`�����:��`��y�̇$�������M�o����a0y�9;��̐	M�~�.y&ĽM�k�DF���(놿��mc�_G��Jr;���x�����dS(��5��*��@���d�"����j{EiU�7X4��$Z��F15�l>�s	�I�U�M�x���>�̱PՁA]L��x�(9�F����|h/�h�Du=Z�:Z5�8�FT���zBk%R~~�cm��/|!eA���Qo��E�	$���p�(Żl��7R+�	_P8%96��4*����K�V����2��N���]Qfg[L�)�z�yǇf�̫�wH�4[Y��1�e'xU��U݈��^:z=����:7=E�l��#JwÊy��AFQ��%��uӱT1��&��]��������>�lC�4ĎKGe�#{�߸�� �F�ѫ���(
b�������տ���0������DXz�@GeV���M�(���lV���Q<(��`�����l	�V���6T�f��������H��4�O3jv�Ʉ���ڑ_�Զ�T(c��h�]}X��J�����G���&\���I˧���ހ����,�q�n �|�T��t�Q�	�G�.��شᬳꕵ�Fm3+�km.m�r@z�Ήl6��f=؏��=�ܖN�e��3���R�=L��GV�p[�������x7C�e�����ij~���3qu�<[�Cn�{u�pn2�ĎajJO�V��~�u��	��c���X���8|�R���4��d�|5���/��ԁW�ի���œ�=���f(�1�vMZ�����$>�!�;3�7�^&x2cq7J]���D&dsvz׶��@<�LT3����J���ϲ{��}(}Վ�~]�0��a�K"�%�1���Pew%=
�*�JK-�E��7qxt�0��<�I�(SbY�7�s���n���\�/���j�Y��'�Y��h׹$3r�_��/X$��D���p�r�XuPVKh5�@.�N�E��kF��1[ÀY�p�8��d�w�?2�)o�C�.���$5LnU%�>��w;�eޔ֩ށC4��V��e�`ѳiX�6�22)�냔���x ���{ݷ�w雿gR�	���%!��S�"*�W�e,�r��0�[��y��|�!�&W��qXt��j?�(�Ŏ�L|�?�p/d�΂�"�sk�,_z8��Ȗ9���Q�mJae�.��=e�˨�a.�RbO*��e�y��ȫ��(L����ͻ{hk.v�(�u=Q�V��6��]��3�h	�ѵ�T~k�2�?���w��Gk���+ޙ����i<�$��Rv��.�g�"���5��&g�A��ާf���;�񲦕z����a�;�����3FV�;��l\7+�2��ຓ�+:1��)Eodx�� Rȸ@��8��T^]����M�n��Tۦ!���PǬ_ԮY����Ux�P �ڴnӯ��^��	�O��%�� MF&WQՓ���Ӛn�e{3����F��Nn�[@���ojĔj����$�P�A=l<��Mf?�6Oxm�jz++7wY�M"g B>�_1����s^A	�T[�s�au^�:j�Dx�92P�p�n'k%�i��B�ʄ�l�;z�Ρ����NJ�ޱҪ��/���S�aTgcI4�� Bv�i�rƤl�M����b��^{Dv��&[��4��N�9��t��F���t4��?xv��Qfm��j/Q��a\B��E�a��젼��}�o+��1ꦢ���aM�U�8�s4D����/9Ym�~�&�eNv��B��3�Q�`e�T��3��SP��V�F�I�6d"��E�A6���
��Uw�p�{D5��!���xUջ��ͩ �6�>]�%�w�ዶ{q�U���5��$��E�Ǻ�I��ѩK�w�H/�����l��hJyE|rX�(�?1AQ�!�jR����\���������'4 �@:����Ե=��a3*�W��������5s�6ϛ��$97��Ȣ��pB�`�iV"��##aqI�޿>��4N�Jv���iφY�D���&�-H$�u1F;����}���6�0�j�*�y�(�`s"[�l�(L��A�?�Ϝ�f
�M�~-6Rܙ�D<�T��þ-� a3Q�츿��޲;��Ӌl�!X���|�.aƸp��݃��/Q�\>�G,َ�@�<C��LcZ3�=~c���M��b��f��O�%��S�TD�j����N}u*�Qϒ�3�������xƬ��̼r^��>"�	�9K���QŝӖI�ݮ4�N���~�
MH����K/��ڔ�B�o������C�.o��Ŝ�B#M�w$�ˊ�#,��uw{�Q-n,�M��@'�}J��0뼰�*�TxG��������D�?i��߇�O2"5����8 ~�PL=��0��	�э���X4x�f�k��W·�W�!�B��1�Q�|���S@����c��U3�(.�{PV����jC����3��4��$e_U ]~�5�ﮚ�G�?;�� �j��y6F:�ïk7��m��w��c���h��Pl����y�lԘ1��Oc��E�m6���	=P�b	H�Hi/��{��p�T����6���#�T:�;����nSA�%5��-Tj�4�1Ŀ#P��<Z�\ 1�%�e�Ch<��-/�3�&��ȚM�g�q﬽j�(���~������4p�i����"�P��T{�/,��R�ߚ��0��������o�-���4u�a�d�9[Ȱ��*A恚0)B�ܚ��D�0y�`������Ғ4^��S<�q􌓔��ͣ�G���[�&&���`��-����!�F�Z�ߗ�4���l��.���X'>bd�XߙǮ�I���.������~���\BQ%a�NN��iʉ�tHy�'�����҂��Yv��I��g%�1%%���$�]��M����
>vw���hIF���4�F��tx��)�����N�0�н���>����#��(w�׸yH���b](x�������a*�v��2{*�J��v��$�q̙����fh`���A��nY�gޙ��N�	�@u��̼4�;6����Cu�~�HȐ��[��y��5Z�����J���K�W ��m�NdY��f�y�+~ &*|��-�`��Y��é�˷\k�|3^O�t]����&*��G�a���|���
�2�'X�u�K��gS�{)E�{&�سb�J�"| ��^w`ɔ�%�"h~c"����c_cPo�LOoMn�lޙ6H�>��Q#�t�vI'ɴ�K�(�:��^�^G��LP��ڔ��{���p��֮��m�
E|t�I�>'�J6�޽�G�S(���VF��l��%����	�L!����#>�h(�	��B:�%��rw�h�1���<�i��HQ�ƿշ_����f���fdd\+�ݯ�1C��Ǩ�੗�3KH$�eY��7v��s�K�*�؞�܋�^S�`f���ú�GMQ�^WgE7|�+��(u��Ҧֻ�X�ϓ�?.L#�\B�lCf� l� �{7&_4��d�[��X� PP�'�ڂ�~iU�K�k45���ʙ粨h^��Y��GDP&V�t �n�{`�����'r�����F�w��A�l��TQDv��y%�[��� ��I)�(��DOW�SH�8�)����O�G�"N�B?���RBYUQٷ��3t�_����u��7�o�T�F��R�S�m�)?���5e'�b/�v�"ƼK	�Q=т�a�P\]���9<�%�`E�q�ͮ\�$���v�l�@�W�4�U:�?��<�:,8˵E�Y*�7���!�3��4^��3X%�	d������u��u�>�U�0�f3��S���,�ғ�1�ޔa��g����j����݁H]��~�3�ФҸV���K�
�?x��2/�FH�����q�����%mw�6�{�g�|z3�T���nk�B}�R�"��=��@�����I[τ!Y-h�KOp�z{�4�qX�]*Z}���ϪqH\�_��T�S�c����`�%ùg�bx�t���#5�Ëd�T1���@~;B_V��BB*�z��\��!����F�g4B��� >Y�(<���P�5F~(�m����ꜢPs� 6I�}D�\�h6m�F	{֜}	���TE��G�l.��!����"���������/�Y�(��r[��t�q R�a6���P_&e�z=�Z������vx����r"��삒.��nx���q��ƥ���k6�xY�u���ķ�%��L���lW��{��$�+�W�P��K'��`+��,X�IC�]݆��m.JE�4;n���F݆rea'kktQ��z�ek ���ݽ�~f�sn��}?���M ��`��1m�F��Ɏ{����H����14>��D�$�SMcx��G�*? �:�1.qT2�Nc;��ִ[=�oGY��`A�<���H��r��(sq�a�y��}��T���9*���[ ��'��g
C0v�(���WjѶ�ӉĨ�Sk\���D��C�7��jB�r��g͏��u��G�M�������u�~M}��UP�3}�k�>�z������9\�Oڃ���fʊ�Q\�:6��5�����3J���6��dӵT,E)<s��9R�U���x֝�K�/'>I��Ĕ_����5t~�k����C�B�҂)}T� ���i؆>��t���OJq�	�q��~�2�����(<wp�	ĘG}��ω�2��qAf�lf��w�'C"X���+|�ؘ�'@���F���M61�����K�A����<Le�V�,��k�����d�~��nq]�D�du�V���g"0O1��Hu4���O��d�~c+:9
��*��-�FTB�� &��a;.,�vc<�KU~��&�������]����7H�:h(�o�T�%�|�:�(?ͯsr&Q
�nP��y��`�H�����H=���)>
ϒÓ#� :Ɓc۞Q�r���+�����D�0����ԛ�q;M�`�zGӀK�����<C�@�jg�;i)���O����^�KB֤|��,�S�?V��7'Z���ؔE��B�UK(�q�$f��#��t��q0�s�9uܑ��{=�:Y�G�̈˝�|ٞ �E��2�����J[�i�&,��6�o�v'SAʐl�!�m����{#`�5w��D0k����#n�At�t�Έ�0�d|k��[C6���q�j"š>qf)a��=�5WHk��^o��s�����iq���"b��ˡ�0��ʭ�LVS���;x{��+�����Ô��|.K�1���q(���r�<��h�|�%��|#�@���@���&��R�P����6�C=yL/�5�I�4�>��{Ƭ��om�O�6���E@����T��异@��4z��U��{~y�3I�
�&�]~H���.>�$�l��}�Hq�����L�Bl��d�M��ܿ�O���ˆl\h��ʾ#l`��5��p�W�2x������;Y
��t�L��!�P�����+K�����u[&��IE�� �����B���[����H����W33S���w}�Wn�;���X��bs&�\B^z���ѫrz��~y�)����]��9���Q�3	B�챭[�bw�����ϤD�,|��OA��.i逪Jj���$$�$kԷ��^�
�S��z�pa�uQ&BB�q:� ܸ;8�����ٕ���7M\��/�p]�3�=��?57�"��e�xFn���)^c�(�d��e0�XO��/�МǵO:��T�O�%$^ע¿��B�$	�a��7��:~ ��@,@4���2������w�����3&�u�Afį[�s�3Y�"z�J���_�ȌZH�if��,�f%�j�tN+��8�xg5��6z�y4`�U��zv�s���^!sg���O�q�J>�+���Ͷ�KChs�bi�v/	pЉ*�~��:K;�b#)E�- r|Rf�,C� ��Z����R������K��[E.a5?p�d��ў�j�N�{������L�飺K��N� ���_7� �6�I�e�G�?�K��e�(�mR	ɤ��n-M![���<���Q�P�E�
�ُ�CD�����9Bi��ni���б�z�y����t���t[��]j�ӡ�&�E��X7f��5�u�/\��7!~�4I�c��G�l�-�/�����V�%hT�r��	ctײ��^��wHQ�Xxǉ��>����1�:',y����Ï
��P_��9������@����C�SVy1vaH�x>Ŗ:?��!o�T�Xǽ��Y���Y��](��ޮ�QV�ćI`R���O����LC]��;~��miF�t�&�l0�f\MݠN�e�8}hX���@�-� �&�{+gM��tm@u�n2��"iΈöL�0y��U9�l��k��c����kei�i��R�W�h�0����8�4]qF���z�����g��7��� ���"��)m��]�".gj7S��Z�U��B�x-�@mb1HRs���ш+ٱ�;3e� a��@�V.To=ֱU��Yq^O�^��?�1��NΰzNm�����4+���`t�O�6���p֘���)7�� �����iN�9�����F���1]��7�e�m@��W$��ԫ`�uB$c�d]�&<`n'�)��� �=�.���н9��g�'f���ﱺ����]�ˊW�6�=�S1p�n��F0.i��݅�A�����:)>�>� ��H6`�Pjw`ާ~;�V�W����K fG6��,l�.G�U����7���/ڞ�֔2G��S&�A8���[��[&�fMG�l�X�m��g'��&d*`��x����8M�;#'��n��e��sB|%QmJr�\ ��������k�EC�,���j]��u{�ǐ�>�?�������>��h�L��na4�"y�Q��aQv^��SfS���b9K��V�J��A'��n�i�Z �K��xW$�d�y��6�s�U��� ܛ�K�Ip��^O�YH�����1��Г��w��y��̠�#������t<��Tq]��>�뇓��"K���3O�%Et�\7S�|ѩ�������f7vK4��{�;&w�kF*R8���Bo�ziJ�š��3�ZӬ���Vo��k��"�� "�Q2�XK�t"XA�i��u3�#�� ����k5	N=搃.ep{�"�.oS�7?���?<�$3�ip��"�Y�.}��#�,ЫN�3�9p0�o�e_4�����=����}N��=��T�
�pM=�aLwzK���qK����+��L!�^U��,{�P�#�4[�C<l��
A��5���N�{����s<4�y9�ߛ�*N5s��*��Ah��@7P
V]��w� 2��^�����ؔ7ȿ�N5�%KQIeKܿ�ъjň�ҭ.�a��[c��N����m����|3��U���Q�t�:^���Q��ʀ����Q��,��Y��M�D���
H��{�i4,-���j�ܤ��q!�o��D�y���M��!��@�*؏ue�K��#<G�g�K�������G`�o%F�v,��h�aQj��W��0r6&�R߀�#��E]��w8#����=FkD �����-�<LA�>��1�����Kz��51�N��˂�D��:��4��8,"�{(���)h���>F�gO�x����'L�C���Q���0��BD��68�*�'_��K���S�۸��V]����ܦ��n�q��N�lį��O�=������\̏��-w�ͷTB҂�L�pu$�$ 7����90�AVI�*�&1M �z�֓���`h�j�H��oޡ$Ƞ��`=�t�L�w(�]�d ��]L�Y��� ̰�DKyڨQt����Wb@a���[��$�iս��H�h��ޗ�|�o������ݟ#t�v�9���oC�O~�.q)��-Fy?)v��8�&M��i�Jۼ�P����]���5j����u��A-����H�I�*s��\�ZT����E[ލ}��4��ǪM�Ⱥ�U�s��$���c�W�� �}����M 魩�w�����H�K�8��a��䭾�[�t9����-�c�7�g0#��/8�$���_�Hѧ��:���]��Į�G5��0.�����(��36�����4��Q�/�`����-�X��b�0r���U^,�"Q��a�������ᥱ�c"����e����<�wb�"���┖���R}�z���|�(
BiZE:_HGx�(�4r^(>N>4�q���z��m�Z[�k��:ڍ ��ź*��ϸ�N���.c^�zp��a2k1B����D"el�7�F�κ��nH3�B�v�:$���6�(H��zi{7Oq5��f~c5$$(Q�|��dgz&�:U'E�yM���A�GQ1�l���?t�?���"Gq��c� ��IK�RU�!��)�!�INDnI7�w&�̮!����ַ����3�I��I:���N�!O�on?]nO���6�����v��y��$��"N.�F�LxE�ɡm)1	"�:��|\�6����D�Q���/1�]fd���'.�0����6I�Jx����N���a�o}L� �Xs	���ÖayFM��}���W�~��pM�*�����"%��{�\?�L�������e�z����L��ȸxp��T)���#M_˨Y D^���3���uf���+ZdZ�'�A�L�RT���η��(R�a<��CY��q�1=�x�-?���w��97�00@��]�Tu9A<1Y,p�D��eU7q����2m�؜�\��4r��"��"D/�Z���Αm������H?��E4�9�9��sO�!�gtS_����&SG2P��5?(�U�6�w�]�L��z+�FP�D~^gAY�N��3�A�!qY'뀈a�L����P�}�k�\*k�>,�$O*�;�����*[D��~��;�T�
�\����a���V�`e�:��\1k�~�z w�65��G?�(U�֢��v�meZ�6�N~��KH�dX���Z�*,���T�()O��0�Uy��N�0���٥L(�\(X�;gH2t�ˠ0'��q�~\#\L��$�ՖS�����>P_>T�����z*��s��'��n�p���Z	�4e�������&�HV��w\�:�������o{�⠟�`������Ո��&�7���C��Y��8��A$���ǃ��]v�P���[qF�=������=#���x\xj��琮�_{ge�i�5��]��ۗ��ِ�C,�h�$I�vп�Vm�8	E�QJ�~.���m)���o���������e��V����:�$aQr�q@�o��j��S�0����D���_���3��8b4�����a/����q�h�y	�����)KEU��gw�V~E5�.0���(�C�zB�M�	��$���q��.꫖Q���	P
)���˓leD�'����揯o����'��oBw�{�@<�:�UQIf�A�/h�I�<Z!��4�=MA�Kʃ9��X�j��T��L����$JqƉ���-�D�J#]U��V{�8:o"rV6n����3���X�vĢ��Y�����L����Tb<^�ѱ�R-��̅��̾kI0��$`�	>�x�0	 �a?�#�P�^����|���84G�g��˕{ ذ]��^8�"SI�2�{�R�Z�&C���lp7�v�s�?ӏ�S��,1�Ş/����y+�������5S�h��(ĥ����/����z�z��`�d'z�C!Ȏ�7������}���un��?��YgDώZ���ǒWV��gwJ���ލ�\0�r+X�Lʊ#�a�N߶�Ef�6�ږwY���z�΂j*=~���V�u˱ǙȚhLM��8�V1��r��r/�[�����j�}Xm��|F%豶�I����l=+�w�Y��љ
�'�A�Xʸ��i�&_UV��*�<<ϔ/?ܡ=|H�_8�a��a5���d�����`03w&��Ek�1O���s�7�~2���\�F]7`Oo�*����fz�� �p,�r�������@���?B�6~=8}U�H��#>��M3�{�E ���{���Ṕ��O��$��Q�Xh��3G�� �A6����=��e;�Z(W�SN���YK�9G��T%������!d��<R�r�/aM���\���o���4�K�'���A�� .��Ǽ��A��?��h8�:�uS��5�K�$���C��FG��ܠ����ER�CO�����SQr�V�u�|<�����$�V��hH��|S��n�x��$�
���O��0�ڬ�\�U�!I�[t��e�µ�!S�ۨ��U��f�u��&f�r��	�N�ݱ)���;�x��rMq���7�s���~'���K�s*X�$*B��\}/���w�f�:���J�tD��� ݔ�<�S��m��/�Wũ&�1j��.ס�o#Wf��nع���ƄBaxmAצfAӦ0�QY�[��9+J�P�f1��X	���$�B�yu]z�}���Y�Y:�T���!��yV�1�yX0�����`�+!���p@��i�5|�Ã���8ޫx53�Ybt�Xo&�"�|d\0�f���
����������<����TB�a�9먡��k��0���Q�֗w���O;26���O���Xj5^Wz"zZ��.D>��/�	�l����Ir����Ah]�g��U[mh.t��@#�_�TX1!�s���hs�ƾ�� 2.��Z
��j�����T�i�qmDMJ-bld��z�������*�Vkv�&4J���a'0�y,�!/�!m Z8��/�\��:�ࠔL��Z�W��झ�:�(���L!�-&���
�/f�H�I3-6������=B�總Z0]��`�t��*�u��HI��A��-����tȆXG����>��X��Q�a>gK�k4��Ϣ*z*sh�1L�q����"{!y�*t����xa�?��'��1��F���O1��gf&���ݤ%��'�ɐ�����̮j���Ǌ�,���Xj_~��.�o��}��0����O��<5��`��j�+1��PMS�K��J��{d������B��U��lWdЉQ:�׽��R]�<~X9�b������an����.��m�	 ��B�P]�$|$̀�2���#s��ö�e��j7�Z���mtN�`��4���B���Q�l�ߤ�O����}��O��gD�*ї��d���P�hP��Ic�)dw��6q9�FG�"�����
GX�������:�g���ш{Y^�o��v��%;yA�ҁG�J�UE��,0�|���ʹO�X�%���>�,Γ���7�a�<��YXFkď��H�?��f����M�p�	�zp$D��p'�^�r�͠��X����$����mnB�LT+���kѤL+��.��"B�ڻ��O��Eo"�lrqb?hig>��Gpc�9�p]n���L��F60mݶ�ƫ}��j����
v��G3m�V��A��U�Us.��})�����A��'������LHثJ��#Y5=E�L<����v�"�&��Zg� ^i�.�����1�L��7�t�Z���/}�3>��̚�JϦ�t�*�����J88�>��\�����c�|��!�g�ܣ�1���c_[z�!r��'|��c2�L�}x�*�������ѷf,I�v��_�ɍ�,��)z���6!��좒�����$��y:ۙ푝I�f@nޮwV��1)%�N�Wi����}
�h/�RރS���΀�h�,xサ��o��@����^:O=;�������c��K�(ֶ�EIdmVur=�����i��������܀��]CcZ�|����˒=q��QУ�ª��T��҉ğ��K�shx�4c��6r��- �ܟ��`���PI�^L����N�́�r|��C C˒�/��G�h�P�{�Ϣ,X3`|�����F��Uu͔���� I�.�X���/Jt:w5q�V�do������f��Zy�1(��)�
A$՞Ĺ<�.s$i�S&k��2"��S5��W+7Es��'np��\����'T>�LM�No_xy����Z�h���(nƍ��4E.��C���8�V 5�������s���#��3��5o�cU��^ǫ��P�1�A��U�5�����UA�V���qr�e� ��0?�=����D����yR�t�x�V����x�0��!:yі����MU���8���b������p��NiDN��[������o
���zT��Ҩ�e���`�	>���
hK^H�'~C6��?��x��s�8�l��k�b.��=V粫�t�mz��ڮ�e�-�㖦+\�ǆA�n���d�.U ��D��@�
w�d�v�HH=AsH�ǲ79���(���+�5��S�1D����&%#D
Jh��~%QX{��X!bL�:l�Z׃>����A�k��n�CxQ,�_��1^�p{QH,Y �6*��:%��TQ����Xx�>�0;��
�17��x=No�7,cy�~ҧ�p�ho��2&�^�'�%�]B���#�������.h�:������6%����Ţ'xo�Yj����GK���M30#O�]�c���35��X�] ��WK�BCU���+�!������|y��aÐ���X�$0�!����h���J0K���LS�;�^��ü�/�]|%/�yW�{���:��&�5�<�3Uh�[Iq��請^o`
ڞ��j	#>�@�~w۰#�~�x��Q��¼��W�E ����1*c��3�#�����;L:c:C%�&�e������/�X�JR� D/�T
w�+�#�:ë�%U���s��y���t�P��y�~�SlI6�Q� ;'*J��ȴo�`��[�jɣ���'��y	�K�����N �T�+��J�ո�G�R��-���
���*�忺��c��=�C�d�	WڻC���}Q��&`�|�8kL�a8<�L���{KQLA�7�
�6� 2cN7�E/@փʎn��	�T1���b+�5r��W��F5���d/�$:���F��6�nڅ����@��7��;��z\f�����_��oP�=W=o$�x�T�W�[���&�T<���Sb�4�����cs�8VgG���	��D��RY��c�FZ�:s9�!z� Y!׹%S^u�U2��{)��I�������|�c��M=�<5(��1�j��w	�v�%-�w�f��z�Rm�H4g��a�W'���k�qK ����<��qF���K7?��PK*Q[-�����{2���[�Ι?�*��OE8��h$�O1�ſ��d#�Pt#��[�VV�B`�V�����#�f�� �[���U�n&�YѲ-�S%�4ۍ!Lg�#ڿMT���\��֭_7�ã���P�7�zh�E����p�o������糿ՆO柆}�6���J����ʷ���b|R�e�j��CVe����v�>o̟t 	���6��tո���ǰ�{	Htג)�����w�8ǿ��r��셹' ������+;[6m+�BT����LY�%�H���Ҳ����Dû��x�Q�	��JD�X�?���}��oG�RPm��^�Ю+����Q�]b)����B.F%
Ѥ��&t����G�A��G�^H�G�n�T[����z0C�`�+V��޹�r�`'r�ԥ�Ú^w��U��m[-Oj��{,������6D�U�N�k�.����m�R��:�.�8�Z�p˦����A���չ��+RC)�zR�7�NE%.��FR�s7(�����"��I��n�s��\��i����!�;pt��HB�����<,�d�Q� ǯs�h&x?|snp��t���������!�L�1FIx�ރ����I|���Eo�W	��;E�r/�'6D`~,�}��ƍ5���t7׋�H��#)�� /@�b��!ټ�h?�~��m$��n��w��_~d6U�A�	L�d�2�v������������e�@|Nd����E��8zUῧB���Dn� ��R ߋ��C��z���[�imT*HL�1�37���L���f&AA��{k=I�7{�*�ױku��c��P�R�S4���B�w-1i;��}���EZJ��-�ۤ[��	��#�>�z�����v��5#/�UT�5
�2�0��Ә���ߜ]Sy��c#
��}(�ے��E3���с�lx�-��%e�$~F���~��P)����Z��?Y�LxOGB�v�E)��'��bn?w��
�]��o�y�� �ig|�1��ѠD=bG�T����"f�|�K�2�{�u�"!�7�đ&P�W�1Ɋ۩-�.}�
7�����m���6�͊7t�<S�A'�t}Eu��8�&+?U?��7��uN5�/��*�HjӲ!$��89��g����O"��Zz�/1
>#m�3{�� �aW8�]���]6�:�!e8f��8�2��6��خ�Cu"�v֦�/Uz�b�pN�X"�	�cF���t���J�09���k��JWQ�M�gT+���ʌ��6T����)өͣc ��� I3���J�n=(]��>�STU�^��M�W+���n���gc��Q3w#S���%�%#C׷������0{���j�h��6%V����i	�	S���AR�n�}��n�({�j�L�z����Ӗl�Z=hQ.��q�R�݋�M��b��f�	�.ΰ]�q#2ʹ ;5v�d,���J/ީ�q��b|I��Z�jK����B_XS%���<��L�e�t����ӷ���D�0X�$[��k����;�~*hWɕ��I�B2jw��i��'�-�R�z������V����I�.	Bhm.v������ �j����S͒����:�������F���@��foA-�0䶅v��FC -�5
k� q�����(4�7���fr��܇��`����c�x�����J�WkP�a
ݛ71��Z�~܌�%��fwW)H�S9q�k?k �~�E��8R!>���	���3�c��t8��Y.]K+'7�/�w;�N�2��? v<�V��]��	�M��Q�[�.#��C�
�n��A,6��0�p+��	iE�3[�7K��m=}�/c�wX��m���v���&F����LG��9���/��Ÿ6Wq�w�����I�n��ǭ�����P]f���4���d�yb,�gKT����K2L��@���f��'ޅ^pY��xN!=�S{�Q��9�"�4����b
�-M{7�)mǗ��ja�K�'*Z���*�i�Ȭ.�S��Lw����2�]������8������$q�S�5��N��xh*����+.i�.�;�wv
-��7���l�|��S�ק��_z�	cg��[�����wy��E{v��@���Lӵ��=	0�>+ޭ�3}2ӯN[��qQ�O�t�y�nսq
����wOd�, ���J��8�_�������4��>�Z�UOT�:�������BV�wj�	�yOO`u�O�+�e�T���+E,�o�A��E����Ί�zny ��Q	G;-���%%Jυd*e/=VP/IT�(�i�"4z���*�� wȵe���z_�&(�ڵ�#�_l�9� 5'B���LA�P��6�k�K��9s�M����3��U��OM�ò�G�?�C�U���`�o��ݰ�:�є���	gk§��]
p�O�*,������K�Bߟ�\�L��wK8W�<���dI��
�f]�.6vZ����D�L��(Yik���e܄�`Ey!��\-��4��)�#�U}'�g?��.9�_A�=�@aF�/Jv�ݚH������B��%Gh��S�kӌ� z�Z��U-3��b�Y �Ti��K%w���L�~?�������n|��XY�a."ob,w��n�{0�yjN�
R�1C��1��掣ga���|���ki�����Ն����HDf��fϘs�'������Γ�w6�2�Ŕ�9Gǘ<�:w�M@/8>����"�~��e��x��K���ߜ�vGOUr�ՉcO��a�Iޕ>+��bd���@R���p2�N��\���̢���f�O�}��6@��22�����{5��	���_>��љ��[S	��xAn��3��7���H�	���_���g���q2��"����$ů~(��	�cu![�!dG�VU!�z�0`���k���m�+dy逎�,/g���/�d]�2��*��:�li̞㐀��=���_��G#�A���bu<&�8������!�]l*�Q��ʩ	!��}��p�MT% Qcw�VJs�J�t$@�m�^wٴ�YH2�I�m�n��@N��۲�q��up8V�3߾泩9� �Srl0����v[��Q�q�s������"}�3���+��5aX�h@��h�^�^�@���,�����S�嚫,p���c��!�a�m::���if��`���n4�Ǩp��q����%���u#���X�$�n� J9 $�(k��ދM,�&��!�I���Y�/����v��}�p�eP������k���]���Qb����K�&gZ@�O@��)$}����\̹�p�̓�)��Kp�����}T��H�[�תf_k��v��`]��
�*3;i��h[��D�4��!h4)m�3H7M�АDU2�E{��
L� �	�=��z`�����RWI�kv�%J��!"TX/eA��{S)��'8�=%s��� ��3k�(c��A�S�����G{>��~B��=X���=`�c��b�3s!�vY�C�#C]�9~�ʓ��~�@���qv�n�Oث�щ��/����k�����Bw���5�p�ߣ�h?Wn7��*���m&�#�l�|��Ŗ0C�F��160��<���Ozq#����!�n'`��9��gx��zvfө�e��C��k=3cb��@Q�o���'���nF��3�z�/�����+М]E��l���jP<?k�J!-���#�wB��O�.�w�o�;��* �9��T��JJT���+���5�����.ͷ���P4����X�����(%����jӘ���x!@����˷��-��+K���g�And]�窵uR�4��
� Q��	+43jȳ؊Ŧ�]��N�o"p��+�=Y�"'B�����H�*�ڼ�1W��^؇i�U�)�F�҃���;uGZ�	����}J�n"
�8nߴ���R6F�� !N��
2�;3���xu������)�L��t��h�8���_|s{�Ku����j�1%efSc�²W!�Q&��	��F��~⢤%�\JUecu�O���Eʘ��&"�+�L���\��É�KY�ى����-�o�SX�r��
9��a^��:kF��gx@�7��\W��w̽�黙��]q�)SMَ�&�].}�=���F�����>4�c֗.���&ӧp��,U;4.�F��|/��0Rr��1]T�-�G����A _�[o=�L�C�Xb l�6�G��t�9`��i�� G��6s��Wc�&u�j�T�(���#��f �Y+8�!�6���..��5W���cC:���9cܩ�
a�߈�o0��.J�P���Ӵ��(��7��p���L��q�	�{(�D��B�k]��� ���F��j�i��{՞�����v��ۢ��a�����k}�Gߛ��&R�Kϭ7}ı
D�f;�����6��8���<����ی���U_�xa�Z^(��F�%;
M������m/��b�d�3�ǒ���������!�	A�	���dh�0R���+U�#,�pYE�m��.�)G6:�UzJ�mm��t�_���~��������,�,���h�X}I}"v� �HSU��{���?��Rs ���F?#O��gΆ�Z�tI��FR^�S���7��I�#�W�y��]-nLY�5�zx������qA�2���&�L���^�],�QР�9.�;��P��g/f-�Q�l���ɟq�}[� ���4T�d�l����[��x�X�s�o�0ӭ��.���ŵ�ߟ���&�Jȳ�|�Z5�=���|7=�Is��:�9C#���R�;lr��ԫ̶R�5�̆;K�Ak�����g�8,��<�#����h����GΛ<����-uLq����2G��ʍ��Gl%~dk�m�Uw���"2�w!��T���0&W��&|��9����n�3�u��������4�����H�l�C��o(C�bw�d�a&�iu�4cp�Zc�~�����''�4���,QYc�X�7��j��;mj�3Ɂ:`��Sj���;�\�S�| �:���'a���(�ĪV���%���4X�)��ځ�C��^Ʉ�z�RT��ѫ3mWdQ��é_y)I����~ż�nK�C�@e��sdn�P�������b�Z}� _�>��;z��V�{0� ݵ6@qQ*H���Pu����M��Cd��Qeu�czΪ]�<�tL���u�|�������4��.!�c�}�8�m���j�+�}����%�CI��_�g�N-�x�}=S�?zH[MFLjn����A��� ��C/���7�c����QH{L�l����SO�D���j�\鑔|��Bb����-;�̖3H幒xP .ܵa�X'5+"�]T���E�������Y�)0Y*���i��v
���y\@|0����%�Ģ�6U��A�XLP��t�f`�#�C�s3M	_�'�:��Vr͐+�� �{�%!p�*J���;�-���@�"[��
��|�H�a��Nsq�S��l���䈟&�Q�`�x�=A7��@Ϫd���18{D%���ո�ɳ���g<�.H��*�����vg����V^j����9�y�,\vb�8���`�Ć��l �����X!MG�� ��g���]��b�
�Nk���g���^	�z�o*&����Z?Ń�����'�vh�r�9�&Jtb�H?�s��ĉ�z�~�!W�{���`O�SAs�]] ��-���� >��Eobv<{)��c`�R���o�j��e�����b�2)����r��f����p/<� �2hX4hE���אe��9��$�����O"�.c��<x���ka@AdNވ�J�Z�>��%�z�&�*����n$:�)WMm��}��DsJG��K. Qԕ�C�vI`����K�4Dԙ��<H���K�^=L�t ]0�o�b~vo���P{�_��Sv��������ב�C֤{�2B�h�&�x�B�v�$�z7�J7K_,��f�
����AD�&��
P�|�~�!|��U"rwP��K䪶xjTV[�}���:�ao=&�"��$Kz�i}C��׸֋ �)�S�J�O����iO��3:�j��7GZT.��D���}�_U�e7��%r�2�ۭ͂�8���Y�^�X�y���g;�'oOn��X�����r���Q��~���M����S�Sl1�K}BZǖ�"��;�N;��X�-UP6�J�fC������lPF����j�P8~-R2,��z'���b�f���-Uy֕~%F/��$?� �'F��-IHth�/�t'~�N��ש��ʚKL�73�`������s�[��6[�C+ۻ�/����� w���'!�q���:��{*�m�'�Z[9b���G�9셈��:e��A�#���[�`�sܝ�$�I�G�RJ�p�9[���6��/�C�{�����
����+�b��d���T�<�H%9>wL�s��;Y�Dp2��S�E��������n���"C&�DF]|w�0��(��}Kt0R�j�u���D�F�Z��)fcYz̸=��_��	��"��\:�@���F�i�/�$a�� ~R����z��<���9(��%���%*��d):����r|��i��2�]g�%�-g����Dv����#���]�uugGA���\�9����@��U�KhQt5�F��$�����\JH �-J��̸)��=��&��xj��ݭ�Z���G���p�>Yj��Q�ܫ�ȏ�/G�n(L���N�'�<Y��Ğ<����e@��$��>��[�� {_u�1	?챑n�N�R�,ኜ,̓cX����$�oV���Xy^=D�B!w�+u�����ɄSK+oJvd��<�i}�(��Y'R�T<�l*�����Y+M�E�������h*��i	� ��hO�{ Tb��yf��!��>�64�ځH/�D��0��c�KIޞ�o��k&��+��� J��r���^)�mn�H�^{����/<��W�y�(xx�l��[��J)d�У����p<�H*-~�$΂o?�zr�o�e�����J�v���/*J&$�̞��u����ۺԝ��]�R6c��n�6/��F�/-�,�d�E����OL>k�EWqDO8$I��]�Wg8l�sg�b��+�"��w��T�g;���e��.�ټ���R+E����\�ż������L�h��`�&��湞��ûKt�8o��?;�f����Bͣ��ˡ���D�y�Кa/�{z�t�u�*r����"l����}����1��M�.n�G?��?'T��o2���Q��q\B��{�_��7�~�\����P��I[%ٌ��{�CLJ�5�x��l�Fh{����[��M��Wl�9�"G�[ڔ
Q�����+�3ܨ��ޤ�����J�l�>b�L����ės�Q9T��&_����r�0/n��b�@'��ͦ\}�����+6(��EC^�?gV�}po�sN	�]|�}ʴX�T�^�/-)tЪ�:���4�:N��O�=��5˥��b�2ʢtL��K�9|G��z^˒�N�'�c4��l��QԎ�����034yO3x�s�8znι#��^n�8��Ü;��[�4w�Y-�V3|X!��u��P�B+8��'�q�7��u��Hs��v�e����x�T�W�3���V�V��R6��*D�JlcW�\i�u�!Ɔ���/p���w*�P���)�
@���[�W��LK�|��C�ހ��V�"��ς��mV�L�'�`�&:�R�?w���=���?㨤��9�^�j+*m�w���>�����u<�do��4	`굃����Q���,w{�,3�J�B��r�5k	�n����L<�W��4䉟5�b@���������%���%Z�+����.\nmHHF2�ʁ{7
BS\��N�n��l���	Vl��T�x�|��H�B����m �p���%`;�(}8`f����]I��׫�q�AA����mw�E��t�|�9��o���YU��K��k�T��r���9;F�h������k�I���kꄔ����?F���Q�6��f�ʉ�6�������$���]�쫩�fu�7��nn�d`-C��'����c>������v**���%��m��� 
o0�G|LE�h=V��&���L�zZ#���l���O!�6�A�/0ݾ,�Q��l��@�����Y�>�%#�]BȲm��
�3UW&��*�D1K�l�}�&����cUD��ae?7 �V����9PO��$��q��������|��'�?y��p�f�����za��3����f}J\����T	 D��-N��4���k�c)�\�w)�F��06̒?�| x�dLsrY>Fg����3Z܌B� g�3
+��� �1/K�i ��ø{�0���]�_=����c�WqvE�#���eE@�`B�����[0q�5��������}�R�w�2B��{��.KV�>5���['�t�%[nwn�:�3���F��)�}�*�ͽ*U4�!�f:���;?\�W��������������U�������[v�3$��n>˷��t��T���AE`���և��f���f��AO��N�b�: &��uIf����O�u�or�k|6!��e��������:�	�u�K�G���@eo���l��Z�4v�����w_Ľ����"�iL:9�b�X�����$�5>D��'j � ���u)6���+˽5y/����t1Y�V�;SpU�u�5�.��S9x/���TU1�)P7D�!���5�8�P���P,
�hMl�yY��=Sna��R5�6�Gq#knTx<y��#�<���L��ݹ�Wjn+e���n���wtuu�\Q��p�[��s|#��Of��U��x���������ޘ��%�R���h0'[�0����,w4�&���h�]�$�W�Q<�4�½�$�r@�r$����s��6�B�c�
_�ok�)�8m"��!�^��{�O��Y:�bp;3{��ެ�׻�Z�3}&�E�2��=#a{0�i���}0���|�A��c��7}�˦2��G١`j�5k�#���7�ε׶�͏{i΂uWT(�eX�P�J>�^m��Ux��˻�q(��
<E|A.W��'�v2�ح�.?�ҩ�_�m��o������e�5x��e��`5{�"ό�J�]������9�_�|�@��Z�~�����x����.�rŽ�R�kg>)����@J����نUasA�^�e��?X��N����K��t!Hۨ��Z��f��u��r&~����v˹��V����mJ�
���r��H�� �T��`Z%Gp`�؉,a/�l�emQ�>�����*x�*�Rd��1��i��p	o9[Te�U��5��q�YA����l��z�M�l����,��wg��;�H8^!�)/�u��/�݁������bN{XQA�ͩ`�0���s�[5���ZԨ��Zh�s)�]7��2i��J��'��d�|Ĵ�b�����1�bnO��;P����
D�)1z�u1R�������ߧ�-��4ԅ�.�uy��E��9��D�I�[�%���9��� ����5H̕���P��[d%�|�+.E�*]v���Te��&Ei��X�Q��J<��Ք'(�� ٝ��?b�����hT�&���٢�ʼ�#N��~x!��SB �>�� �aWwkQtqϬ�3��j��+lQ�]�R��Uy�i�sU'�Ta���l�������p�<JG��h*H�>�B,aE�a��6}֍���Z��#2t��vA�L�ʙ���������nu�l��)�0����ٻEOл;�k�gR��A��c�����O�ං�7���sC|����o�4���֥��D��$alt�ۆ(�\Fj�
͵�9�M����ͻԾ!6x׃[�Jas[Q��YLx)@ �����;Wo���l��~)���&N�g�{Fo�f���7��Q45i���Y�W��Ŝ�6�1�'\Q�L&zb��k�y%p!T�����a�	���xb1���У�-]n���t�� �ľ1�܋~��=`U� �rX�n8@�����#���%�q-���vi0�$Z��b3���h����	�i�FBo����J5b!_��W��NS<���<˵��iL�W��d���΢G�'�4�T5w3Od oU�te���r���]�?�vtM��O�
��N����+o�23 !a��΁�0"G���
2G�k�W�sD�x�*��,a릥���7�7F�����'�3�?�Y�cѭ���#���T��I�M��6/Ж2I���u��Og�?:�@`K��fE��v���'#�b��(�3����У���0`k�]ҫ�ߢΐ���a�n�I�)5_�ބ�(ƌ:�r�L�K�c6��'���Z8�`X2׺��*�\��:]f��뇊F\!2�V�����ԣg�h��N��%)m��X�J���e�>6(1L��:`��tn�a�GZ\�L���sٍgo�dcH���_�45ـ��E��h$u�"l�q�D8��_X��S�ؒ�0nQ�MQ�\%��� ����p;Ī `!��H\oB��7ZȻ�����ά_��O�ا?vE^��=!�pO����U`(�D�j���b�>�����i�t�+�A�G(���%M�{�蠓B;��9��U��k�m��k,����o���f�2y7���gߝ/ y�0>
Hv�ڻC�֬ j�}��=N[f�$r_ÐB�Oe��x��;�#[<��=?H��0�<X{����[Q�W��f�'��&ا�79<X�b9;�Ȭ�yW���m�f:d���by"���i���d�j��D�nnYʫ¤/�0GwnQ\3�� ��!��}w`��\�y�̛"ӱ{W���ŮS#I��7���R���Ӡ�1ʤ�o-���j�ӎo�l"�˩���۰ve�#�D���Xy�ЗXT�FЫ�C؇�����w���;�1��Z�Qzh�K���؀�ǢP෾lD�����qM���Uy�� ��"Ӓ���H�$����t���-悽��RA�C�&�0�'�1�B�"�Xyjw.�Q�PUY�6A��ꯓ����E�?�t�+�U�z)��3��.�2�I���p���q��#]���Ncp=��`��V]���ys$e�T�O���	>�o����&�ES;?���Ǧ�O|	T�om-}���w(���rHx&=��i}>��Z��Q���ċi?��R����`��u�V�ف��^&�N�
]��]��^���)�ד�����1����M�5���BS.x�h��d��Ig��l�ɢ�w�N�W=i�����>��X�W?<6.�Ҁǐ'��{�%�+݃V	�v�|�8EQ�Vo�ʁTr:|�f��%��3-���IT�[f}y��:z\�O�S����'ù���P!]4��ѣ��X����c���N�G�i"9Xx47�Q;rNC��q��<�T�(�T��h���\+�B9����%�]��.�@��j}
�M���[�'�~h�X.�m3R9m�`O)N-�����v#L��@��c���aH3k0�BO�YA�ܞAA2��#���_X���_� `P1*�f'�$��֑����A������K�O$��J�)��ҭF&[�Rq�1*���C�e��ȜNg��V�y��YV�2f��+`o��G��O��?�N���^�J(Gc�������J�a�[�'��ȴ x�N���7���d=sQ�*�b��j��
��E-�6z{@���7t��*V#r(�py��tf��|x��s�}^�~~]��j�5j�\*�&`[as9�r�Z>���}����G8#��T�OU���|��O�	���ή�P,�56˥组4y���y{5J�C�L�W(�W�%�'pHV����yʇ�h+���>�86,�ݰ�����{�]�Wb/K#2v/�X�ٲ�DϽ*pkj�:�o=�6�cb�VN=F�Of��A�!��"���R7��ż�k�/����n1`�����"FP�sN�8�~U�95��A��i5lxt!�,?�|��O����"����ƢS��u��#�"W����H}L�ϸ��ԥA��p�1٢'��$�J�I'3]���˨�>?#y�y*a��/7�*��GFӄ3�k��-�F��;��b��bֹ�RᎪ&�O��s��޳�(@�t��٤�D&ы
ds��	>���|�-�p�p��]�"�d�mB�7�MGN�r밮M��B>qôD*�l#�����˘-ɡ�f�n7��%]�|a�P�`��_��Sr�d���p��S�m�������X�d������4�����o#��~�z���̱�-E����id�WoY(]j[�pEp��[��I(f��`ʈ�Љ0ΝB|(�}����Q��v3`~iX_�9���Wd.ǙfK�a��|�.�-Ix�{6�
Ԛ��΁8�����E-�xkx�x�ۻ4_������x�m�G�$<-퓣��ޯ�^Z�T��R�d�#�ei���6����|(A����Fe�H�dDE����v�z�w���w$�Q�M�L�b 	'O��S��.f?C8���,~d�"�R��DY҇VS�s�����3��I�腹�rwƃ=�h� a6���2 �K/�M�S�`�����.�$��Tco�0 �,��f�$t�%>�[{hmB.rȞ�4>�f��-Hⓤ���B�ԅ{��� dSGh�<Î�� �',�����~��hA�zz~~jMߣZ�^���r��~xwk�]���䅒�ۉD�\M�P���$�e��L����ۭ(J:.��"�I�Z$��TծG=�n�u��n�J���s7�\��s8ug�<p�tu��U��B޻{=Wyٕ��-z�̳�}fŠQ4VX�m�䭓�^�/H9t0M�<�Ъ2	*�a�Oۦ�X�T'>�u�(�?_�.�G���tw(�^����Ù�i�ԕ����R�+\"jl %���!���L���w�p
d����[�[K�}���Rl&�ClR���K���ㆲ� �xW~�^�Q�x-��n��6�{�NgS�/�r������E��j��䘺?�Ь5�njU��>�T�:i���La��ib�N���Xx9Ԫ���툷z�����K9����.�w�s�0ڃ���C�o��Փz��KӿG@�X
�ܽ�U����)�K���C��lT���׫R\�Wg(	�,r�����vQ<�=�}z�:�\uH�cYe̷:��]�[�u~��O��7p��M�!ᗎQ
�`�����5@�1���s����HJ=��61�1�$qO��K����m�Fh��НvO��d����3�����<%:Vg�3d�1!H�����D���8ē��^�R��{/�����+EQa�,���HP
�.C���0����gx�&3_Ok���uo����?+�u���	�K�
ވޏ���;�l$�Qj�|:�0�rݷ��T��mn뢱��uі���)Rd��OX�ٿ�\�q٥�ب��`_���_5Y_�^�&��~uG������H�^}LUd��'��n�%�e,wd��x)�ѯ�7Y�C��'Ș6�暲��n�L�n�q�W%"��$	���T��r�6$�⨕�-�iԍ��,r�&g
+׋�7�V|���#d�M~�3Z"�r���$��g���NP./ѩ�\=7�����76��w#�݂��.2�0ՊٞP��+9{:|I�~}x݆w$��E�zԊR!����.A]#��r�G��sQ$���`��Nn��t�]�v8�k�,�$�~�֚�����S��n$�Z�UM�#^6���H��"���͢�G�t|�I�>��S��Ά�7S1ZrUC�X�wL�?��#��$Q|�4�4�}=��L��+Qc4] �h�ۈ�`[��7�|�A�M (��Aὸt�/��f��L�NLl�+���=oIS,6U�Lf�fN��3CV�����Ck�&�5��`�]܁�)�����$��v��)��)
o��r�������o����K.�&� ��F�eq��K�T�_��޻Q�j@Ň���h�y�M�F�0:xE2R4Ч˸�̦V����!���!�^H��ʓ�:�ۢ#��	�Y1�E��fW�l������W/y�p|Bj�&rټz�\މ��E�!B��c���E4q?���A�|m�`��=�;��ʼ�	��3��;��3��1�]CeI��$k��m��ɴ�E��c�����.�� e��������÷&�/Y*P%�7������g����&-�KȩS�%j�J���|�쫆)��v'P��f�/ � z�ޛ�F[�hZ��\^\�ޢ@0�\��I2��{_y�6_�4D�2��`V#���<��`j��ϡ4���v�2FG������e��t(/H+,��� n~O��	�!��a<�(��K��B]��T�����q����#��|��G���2�]�H���X�r�������Ğ]7�Lh;���Is%ŏ���b��[[�|�!�9(D�hZ9Ep�7�~��ϗ�����ABkZ+6[��S�t]q��p���b�(�b�K�VE�7�B�����Jv����"2��Y��r���@Շ�ͦ����0�r�7f�j��P���=���`$���2k~	!�aĪ���ph��K'Wƿ���&cƬ���Xa��sL�_[�ô_�$|T9��*'��s�)���A�rİE���vfwYt��:ߩN�TKni���ӋܓNAh��B7D/�y2�@1�x�V�ׇ����;�K�׫��i��f�=P]l�SS>�m%�����ӝ�5�s׷�B~G��u'�R�`�d�0��SH�t�s	�a�x�b�����R�sR�;s ���{�`OZz!�����x)H=�����]\*�y�3��`WGӸ�H���&��%Sx[6zq)��x�=�i#�����s�i����E|H���p�.���FD+{jbě����N����2RNpQ��6i�a\u��56���W�nn���
��(ܸN��b�qt�nI$?6'y�}�ѩ(�?4�Q��H�l��3�A������T�%<8��Uq~~�&���:�E_���^�8?^��ޚY���G[���K/-���h��)�S3H'yK��!��+c��;�sI.5���#������ܚa5[%�L��vj�AGEC�
+��⁕X��1��H��B���������y��{��q�>+Xx7WD�}OӢn�u�k@�EfF���{b-H�Yn�fR����ћJ���o�g�jt�ܩ6��%��G�Zi�q�eGڲW�\o��X��{�J��E?.�Jf�|t�sA㧂S���6C&F��$��ȭ&p���~��!]�]�p9)���%�,���?��g"�@3�,�ġMAw��1�V\9���"	����Q=O�������`(��q���EG��s@Y>� ə�t}o>��񯎨��+��*�c9�Hn���qXm[wD�J����_�J���H���3�`/�^(h?����?٫W{7��N�@H8y��x*�Z8���)&*�66r�d
�tcFG����a�DRb�!�5����xa�?u�u�If�X0�&��$�z��P�]�^��ُ^�	��Z����<����LjC��}�~���R�}���W�l�Jr�Q���S7��P�Y#�t0v���b8#[�6 ���(s�Df��%;��qx	1��z�jsj�W�T�9%��x��܈п��p���ȩ�E_��O�����"��D�td=�`SwL� !�Owfޔq����	 ��{��G3�����U6:M��"��U�53�y��FZ�����x��q�{�:Y����H�Qv�U��2�J%:��-8������!CS�#&���J|1�°�	�=0-�.}���,Bg>�|*说�\?$v�V\<�..fL:��K��|Y�m6�`�c}"��uw�Tɾ=s�߆
1+���b��,=ŏ{�21�0�f?������e֟����迌!����g|��������	�n�"�=��`����NL���մ&5
�q�A�����"47R��n):�N���e1�`_�޽�����q?l_��VFTW�*+�:�Fq��E^����zτ�	��p��/+���ŷ0xK�D��/^���@|˾#�=��v"��!d�J�>h��L_ŰΨ�Y����gˌґ���$X~��f��P�:⹝���$:��x�KۥM�FkN�ܥ�K(⪪	nj%)/���,ƍ%U��)���Mx�C+�͓�都!�ˇ]��T�!�4y�6?�>��)*v�ȑ��Y��f�d8�l��\~KѤD_�k;�����]��CG�S9�A���;p�m�,�� �>�dM��+z���j)(�Du����%aI�nK�O�N��sv�D�e�?S%��M�5ǥLϡ6�K{�/O���I�FQ�4��TF�%��Rr��X�7�ea�O.X�%�74�76e��k�A���!�8ӕ/y�3YGe���5�^��yk�:P8L�8ֺ�BW�"�k?'5�G�E���3!��B-;��WU���s�Kt���B�������F3���O�Q�����a��bS��":����W���b�� K�Ž%�w�3�I�҄1�<��Y��^&Q��ѯ�Q��(>���I� v�1T����9�Ru���b ���X�傤��l��bډ�{����j�X|5�J	��7x�}���	7�!��͕;�r|0�~�:�I�`�ݬ��3���!�ccK�%�\���`I+����2�ZpN/
c�CQ�V��^	|�C���7`�����(�O����)^^��9{�+Կ�`;0z�l�*6q�����9�����S��-�]5�5�4w�tąe��'���5�3�������_*���5a�jE���D��k��򪜍$?Jby��n�kY����>���2�lS���s�6���~��d��o T�#k
�ޠɉ�T�����s��dj�zy�����%al��<��gcR�T�5��N���a�����7Q�kH�-se�ʕ$u���*t����^���~rS���[ݿl�t6%��T��$s�������m���<#�x����Q(�5�?@���6Н(����z� ��ì�(j��o=Z���R}ĺ#}�^:�9E�,r�� g�u�#l����59 j��Ox���by �,��?�!�I�Jm֝��`#�h�;}���Eb�1�F�\�u:�qx��pbiL{4����bs�똸�Β�~*+� �9�7,
1���I5�ܥ�\�ٸ���-��K���RP4MKJ�w��I���w�6ז��	�W�jt?Q�4�}� 4�юS�[B5�QáOM�l�X+k�qw-<�NW���c��LJ���X(s��?�YJT.�{Pg+�]������f+R�Դ96���-�����X��u���;0�"����=��<��N��./fR��� ����^i 5�h��~��*�ڋ���eQGM�T��g�_�Ѐ���Ȓ�o��Ρlij68�}=Ps�e��v���!���k9�<�,{w���	t68���.)X ��|��7f��3`]��@|���2�`1+�����#%����j�6��P�Y�V�o.ᷕ�t�@��<?�[�H�����{�v�>r���)�G���+�aa����W�X��L���y9� l�z����q�[�ǠB;������O���ŻpXs�[�_C����N�~����e>��e�ޓ�?(�ʝ(��s`��O��Y��� �P�߅q�X2If�z���J�>:�Ǭo(E�\L�(��Y���!Glϒ�+�?[k���9��K� D�@��t:�q��o�M߀�kPQ6�;0@�W�m�%k���Ű���O��J��;Y"L��(���������i�M&�q3Sf[Z�}�0�Ԗ���e��M):ˤ�$r�X�c�ф9�)��[ɞ��ˈ�!v��c��$�L@`dIj�
A�=��6�+\� �����t�a���tE'�V?O�q)��W��XB�4�F"��]3�h���{bpԋ��u���&.�lm'�m�xi���,T���66
�^Q����t`�d�ݔ����,�F���G��u!�}a��Z���h���TX�F�����)].C9�_��=rԘu6��:�3<��
8`8(N@��zR�����?CYb�BU����4��3t`���c�C����n@a��D���n�ć��t����o9�)��s;�^��Y*�.���<�*��TD@O�?\��/�0D��U�`¸���c��ݣ��Ў�K=+�(j�78��P�R�$w�f��Wxߗ_H3��C/�����f"b�Y����Z�5����ە)���KL��)hOz)Q[�6��|>}tٗ_�[����UB�B��M�Wse��#s`]�n�~q��;p.+���݌���� E�g�G��c�En֕rG�Ӹ|��&���?�v'���hm��s�/��S_��2���ȼ�c�HŴ������	�b� ^���R}��Ut�8�D��'�i���]������{��΀���"
8u_v�D���W��h�O�n���!���|���0"y�����ͺ�E}8bs�2Uɹ�������6�]d�ϕ߂]���z�w5���f�8WO	�?�*���$��x��H�>�4���و_�0б���^%c�@����}������u�_O��9Ef�1��Y̶g��Y!K����6&��lI5GQ��c<qaߜ�+~aV��6z���I9����r_O��j�=�kEBa�� n+z��
��_��q�e�`�ݯ���X��r'�bY�v�w͎^��U|
X�5f�G%=�}.Γ3�(�x��}h��O���1N;�ۭ�'��3�5�?��yT��:��6�鎑l���� �5[T`��{�?�I����;�����f͘*��y�]�uj�+�����6bT3�_���)��Ӵ5��6�����i�*bpPin�q6�X)�B����,D�%�yJFz�����QT�2�&OS	Ǥ�_hNo8��GVi�*U5��)M�؛��swq_��a$2P�Q���%-�P�"��$�!-��ί����k�'����]���c:y�oE�]QN���$��ٜ<ד�GE��'��z�N��Y�m�d���c��F��R���V��t'渡�ߡr�FW����a��ku�{72�RI ֟c����[����_2H.�#K�s:(d��N�|�X��Z����dGcc%��$����WyM�_!�R�e��	�@t�ƿ#ͫv}=��;�k�7�ZxjMTm��^�eid1��E`��b�S<���"!�����48`%����B�8FV��&��'p���	_�I�z�H���>(�$�� M�u���En��[>��$l�
��]̮R�/]b�r@��'�
�.��qK�sŴ�ܲ~6�wt����V�`ee�����]�8�T�H���ͭ��wgb���_�ӎ2%��j���}h{
#M|J"1z{Fl\SXf��0�b@X�l�L��5���a
<���gw�]C��ɉX���z�i-�-���|�2�Ǩ��˵��oe�,�%_�6f���բ��qj��q磠"���k�w��#�u1���N]c��5De �u
�`��U�7��L��MQ����>9&t>���ֈ��8��4^ud�_7:�P��J�T��<��Bff��:�����O��G-��2�/Ň��P�w^�`�	(��:�|�"��C���E;!47C�)�2!�J�Cd�@ � �.R���o��'9� D��^d��PЪysc���RoR�v��fh�H���;�\��S�_MC��r���2�$2"��c��]OI����{��a����:}�L6o̄˺M������ ��|M�[����KIa��7MU|�ɥ8�(aq�`5\@2�<l��P����_&FҾ��ϥ�3���<�||w�9�<�[��Q����QT8J��/,��-hI�I:Dl�R�<*��^a� �����Blƅ�ו%�d3�-,�E�/�灲MV[����e�S+�H/u���® ���;���"�3��ը�%a�,:&��_ڈ~or��S����zLge��};NҀ�4�y�=�y_F�=B�5��#��طN��w��/3���9b:���s��xT!��Z�(�W$&����{w��iG�|����qQT�
B;�+�n�D-��_x?}g�5q�H�WV�T�g��D�ɭ����%��J��i���@�x�ii��st'P�!L����)e���;B�X���ۓ�
׾��s2���D������r2��#�o�Q�K0�!���c����3���5�~����m!�?�FF�����Bwk,�щ`����V�o�?��Hp-���7�
�rU�B�� ȋ�W��g@�k�h^2��-�X`ڻܝ'�}	!���JQgW�N�M ڞ�)'���J"�Z+���_z�No��m���vEY��{*�X� y��=q0Í�w f�/��糧ߝ�jO���x#h��F��#�x�q�iԨ�{vBO��g��>���l6�!䋗$�/5ř��g62߁ ���q�z��W�Iߔ� �d�'+���P������ ���Ӳ4�H�L�����9�X��-��u7���	�P�>5Ao���V�TX��=�@�؀!G�~/`'�0��\L�MP�έ�v�5v0=�y�ZR?�Sw�q�%�R��X�k�*�Z����?r����+�)������`az5)�s��l�#�e̹]�����%�D��(,���h�8Dܳ�1�
�%�Ep�G.�'�~c����Flcәt��Y;�9NŜ�9U��o�o�iY& ?�J�
re�Jx��n�<-`�Y�=�s���9Ay��eƏ��'�" �Y6c�X�ekv��T�#g��#�5�5�	;|a�za��o�M�f�Nt�h�Y^��֒)?c�͆_��	ͯ�Qs�� �S,��J�8Ts��/�g��V����H� �-�ؗ�}��ߩδ4Yuʧ��0�u�չ���S��o��^Q�z1�u�E֘��ܠ�"�W�;��K#���N3OU���0a���K~��Y98�w�.�;���1�:�ݣ�r�挕=Q9�m��D���~=ۛn�N��DmWbm����Ҫ���ٙ��}#��� 'g���joY��<U��.�3������/'�a��?�Ȳ�@7]gαp���b�ҷ��@\���͖��sH�I~#r�1W��x�Y�����2�2�$$B���X6�и,/��OAA���|�;�G��l3�=��8T�.bshLM�Is KI3\mᏴ<K��
!5yܛ+�c����0g���>j��"��\�LQ����Wy�R�;�,VIG�#�F��U�� YQ�����(V0DL(/�8U����*�VR�K�y��;hE�T ���*�����.W��+�(��Y
�T�����Y�?�~�k.|4O6�j�nۛFͰ�v��DN�Q:���[�{շ[�a�g�Q%l[02"ݥ�r6��V�sM���?>.�� ���%����׼�#�D����d���t����U���K\sɁ��91���ߔ��1���v�]'-��������ٺ̕���I�g�X�c�#�c��[�7ԔH�Ėy@�騻�e��/JP��:��0��$f������k�R��J_�h���a	��v��pN�P=0S�'[
�Ǩz����P`B^p��c�l9O��A!Z�P�wL��C��jId� �V�����5`ڗ�,M�K9���x>���l�����zܶ�����<3is�MMu}�9R?����?G��Q�?5��S��z�n��^���5��Y���D�Xj��|a�ɝ�~e�-�rԨg����-	�HĀ����ͳ5���" $t!��(3j���G�

*]�;y#���#U���f��.��ȡ�����
�I�Vjr�5v쫯��*�;�ѻ���?�lb.�a��I���?��$��XEW�b�����kN�Mܧ�Q�^{F��������۳R�b���FB89\���}�����ޣN��$b�!���`�Asxʰ%��6G�)��ť�.
z@ȫ㠨J�ێ�v�Aw~�f(��R�{�U�+��z\���L�J�����qM`b�������ԏ���AݡY �`��T��ΌjB���e�N�%}h�e����F"��=��Lr,�]��{�	W=����+C˦�n�y`Hp��d�D:$wf��|��]�'�$���L���  ~��k��M���/��Cj�Oƴ�k�ۥ�<�^�t�"�+;rb�,`�� Q��c�"t�C����<����j�"�90���؀�@��(�ix(�f���r~n!c��c�[d���e,i0mq(r��ȸi�L�sڲ��8k-އ�|�?l�Ԕ��K-�����5�-;vdA::F�B7GzbTH��L��������7N�����$���	�ƶvwO�(k.��K�@��p�l=3s�Ӻ�/�A3.�S71�WG�ԓDV_�
��Ĝ�E[g M���K㼭M�Ğt8�s�ޠd�8Vv@�려r���"o�׳vg�5޴R����>�N�*>�5��g��1���7�m� �9��B�-��r��,�����(���[0�/�<�
���W���k��>�� :5r�X�m����/��?�56H-W)2Z�!�[}��H"LD��U�1n� \=w�#�b�M@�}�/�k�J�:���
��,&��t��wzhҩ�g��r�KG���i[�kl���!�7�[D�����B� |L��AQ���r9;�������s�(Lz?ڇ�N>׳4^�5��wpȨ�Z�[�{�P����o��(��\�(I��;�i����n������k�!�k@�6�aSg%t�i�=�ia���k/�!e��&֝�w�p-��4���0J���֛z�,�m6®agk1�d	���d����lZ��(1C֊��\�a	�FJ
!%\��_�f�76˰n#fС��8ݜ5__f@F�x��'Ӯ\�>}�+�C �Pyeb|��i��ſ�~�����%h�;�9H�@�}6��?��Y6�����p˒�%�e�"(�f$�
a�dVCEvA|$���ߣ.8H2�����!`�F�a�ŭ �j�w����,-y	�2AcB�	�T<V��q[Dਗ਼��>x?�eU��A��2)t�l=�W��щ=�8���^��L�?��"=�Yvơv~���[� �]#��2���ĕN�K���re�)�=ˆ�u\�{\]/oY������l/e�XȰk�>7����T_jMr�@�f�����c'B,�6���<e� l}�IApZ��}�����c罘�^D�<����J�n�i�Vi�"�X�����<t>��ߵ��0Qf���<Q��w�h=U+qo�����o�b)B(���&�{��E�F���#vZ�R�fj&��Y���b�<mY(���<�*��ݥ`,{z!מ �r�((�[���w
f����|�0���܆)_�) �x��u15�$�wu�%:_< .��Э9	���b�����
1�k��6��;�ƾ�˃]�{�4�qH��;D�p7"`��eC�Wߚ���f�i���{���z@����:E�o�3�=���@k��Rw��5�4� 7�el�{V=jW�
ߤ����'�"inF+�Q�/�D�����{h3�(�w�@��>�P��{]:�V�ع��ً��D��`Ϲ�qO]�Λ�/�k%t���o^�T�O�i��)�&�����^a����S�cr�K��\	���kѳL��~��j
� %�4����{��V��6��l�J��Z_랼L��H?���U�+���;��1�zL��Oe=7lD����C�7�����Ũ`&��ʸ��q��PMx�L�q)��A���dW�.��M�
��U�g���g�8dv���$5��LEp��:D9�A3P��,�S����޲��'8���%�ZD|]��P��i׈hh��
DQ(A�.��KW�j��e����a���KY�u��q4�VRۺ��p�s�;���(=2����\��0�jW_�|=z��N���My1=�,�d�\3�L W��r�#!TA�^�N�]���zu�Umh֐O�a5߸N%q���t�Ŕt.x�G
9��n�꼷T	�G��!pB����^} ��; ����3�c��n�j�!L��h��5p��{W2Ȥ�� ���Ͱ����l��Sr��)m|�Щ�&-�����b\=DPn���H|>���V�����b��.�-�k����qj؄��9ʻi��e��3l���'���֞�'��@��:%�.��3D׃@�7!i��&��o��qvm�2	�X\��zĉ�PU>c�En^��j�}gX mاN�O��cqχn]+�=�Ɲ�������^�l���a���{��ha}���n����KH�|��3����^����l� A��C^�#R'�5,�k��c����H2<����_�U�PMEa�F�ڸ��ԡ�`�	�|��ۮkլ.�q�V8��_U������	�C��Q.��Ƈ���5�mⳛ��_�AA����(c�'A�qFx��O��DP�z]E��J�����ЫF���u��_6�P��:c�g��@��Ír�9��&�Մ ����:��~!�5������"j��%)�,`�4\��L̷��+ì�ږh������_�<�9��|��d��:b0��Y�lM�L{����vd��"A(B~�W	rϬ�IL��(¤l�ԓ�Ҩ.Q��A,���kYp��ج��C�j ll�F��_��K��������I[�l"tԖ��Lv&����^��-ɾ3r�M�{l�*�B�6����T���Ӏ�ۑ[�z|XZB�����w�(׏z�*��j�z+ũv�j�%��3�~�:g{�j@eD��=)��;i�>�l��,i,�E[����ȧM1�vhrv�����/���(�^���a��e���x�}���&��e�v�Ȇe��!���I�x��$Y���|iZ:x�����8�ܺ� �Y���&d�_]��$�k3z� ��U:d�/�f�9�^`)��$.f&Q�3�A���;�������^',x �|�Rb(��} ���w�F��[��I�}���ڣ}�h�|'�.��A9�7��J0/�-�0/� w��[Ze�<�M���0�az�כ������e��5���F7e�2�93͘-��[�?"h ��[�o���8�S�c{M;=�҄��z��z~)%@?���8�}9�kA��@k�m5�/�*v~݃<x|��曑��9fQ@cE�.eH�c�,���u������Ks���dx���$u��Y2txÞkH��t�U���8Yg`��5`�ٌ��CY� �XM�i�����-1@��97�9�����}۞s����+�n�0���j{�s11��dPL$1����[~����#iOo'9��n��N��Z�8T��u�t�U?�읽�����4��CZ������=P���:������!�����.J�{�������$�AJ���|Ea{O�&�;�֌:�_��ͳ�5U��������q �s��6c��U0ސ^s�������ɁRӵ@λ�7�����l��=`WC���\^U����E>!>]a/��Q��y�Q�����s��!�t�+y3�*x䟡��׼l�˿���Eul}[�G�=uj�h�B<����2^X��?/�?����Q_��3������`v�"E>&pZ!z��q���B�(-{*�JX�\�-5+�u{�R}^ZAS�dML���I��/a?�*o#�q�Vl�4!J�}.э��G5�&r���<���g���޺�JV�	�ox/�����wK`�ENU2ǂp��WA�PF�z�ݝ�c����п/m�U<�m�Ë�_Yj���(�>�^��w��(���bN]����2 B!yyæ_t����H)���w��1T��mk���a�Q(�i�(5Y�4�
�f����'N|��O��w��{�y���i�~��I���m��P��4" _�t�;��PHuaba��'�@�rŏ�(W
Z��1J"H���E}J����Q�4Ă����[��zs��x��D�^m�\vo��G@Ѕ' 0�<����&���r&�s�B�8��B�q�]�G���v�b���}���M�Bc�������GfJ���v��/U���O~Q���.����������۟l�<P�\�	6Ȝ�k����T�\`{#L�֐�d�&�I�S����R-l+4�b)�1�2�Jcd*n���	���rα��5�`g��C�#Z	� ��#7��g�������B���Vo�� `f�kK�e<��*a�oCܷ�@R)�u��Gk�J65�p�Rq�đ	d�M�6����ۨ���W�� �b�n����KÖ��WG���9���H�F�{�8u%B�y�o��al�^Z±^����^O��ڀ_R]e	�M��ó��1�QWlLKK��Z������6'1��04?�֫^S7�K�̪yD�Ȅ�xZ�Te��o��B�&r�_[<�A=��|��� oG`�U��W�I�i~�<��R��� ()l��zT�T	����H�x�Z�\�݀�_��4�j������d
�����W$�@�w+R�[J��+˥Q(u]����}v�@��:e֤��� ���a��!A��O����?奤R�¨��&�j��I%F:yb[,�j%�AY~�P�s̴8��`/M�C�`ī�܄�ϱ���I����.Q�bO-�v,,��y�e�;�S4x�L�^�(;4��d��Ud�Rbd5�����md�|�GᚥM_�����V��0_���,�ղ�a�����c�(9�у��4�"(Y�&�m��w
+��AD=��s�ww!�)��P��U�e~���â�S���w�IZ���S.]���&�5�|�M�o�����)��Z����8;�.V�)7P,E��
Ȋ��)3Ӯ��V��ҵ�d�۽��y
ǖ��J7��	-J�&�e6ψDò�[��?��~���f�M�)[�؉��Ҋ�|�7x[CA�Ub6i�,&?��6K��Qli[uQ͎}1�1C��(^����N�t�z�+��㹺�����Os6��:����z8��%�>3W^�ue�m�\������Wb^6��İ׹�S�㭈�#!L�,p3w��:F��4�|	��
J2� L�PX*.��c�e��a9�k��5�t�dF��tQ[6 ���՞�@�$�B5��/ti���m��9���M	���`�ȏ�܎&n�b`��K��x�q���I,:n�������B�j�#Yc���-w9�2�#(e;{����o��j���\#;"�D�h��&.�#݉
����9İ��wn��"R�A?|���*��2u3���5�@!�,RW��BQ���1���{�J��7�f��_�RP&G]�+�vq�o>1�;�(��=�I�Y��+�r,�LSOw6wn!�`��;����P9݈(�_d��u��+r�l�[��H�:�� d�W@�ˁ>�PB�ħQ5nv��6a5/�5L��z�q��y0�)8�'���)r��������M3�G�@>&\#������p(�f{4�Z�Tu��N���;�S� \H��~i��Xn��5.RL���v���@���g����W�K�+���msЯ֑��C�Ă?��F��6��ym���-}N4i;��_����1�M���Զԕr���s�OR��cU꯵��!��I!�{½�{����M= 3�!,����np���f��1 �J��8�k9QUO��$��'��� 4��<I�e,\�r��?���BD6�� MYJOƦIה�L���C��?]y�,?p�ZM������ �o�CUڶÑ�<�q���̤�{B1�]^����}Qg߾�?Ō����t��(���x�zx�6�S�mL���҂.�����F��S�aܼ�K���G_T�k�~}#�xe
�x���i�q��"��O%`�ګ��đ�z�#T1��sW���@��]�3h\�o$�_�<4s���e4����~Z`[�8��PH֣A�<B�HG.�x�bW�>��4
�`5�����vՔ�����p�jQ ���<�y��p��I��\xX'Fbo� ��关Y�2J�7r��J��'����)����v�ϑ"�Hۥ���\�����P��/ky�J�[����C�?����9y� �@Y�Y��>��Tա��-Aˬ#!E���>/O/����Z�����^Ն�5x�`� g�)���&����f�#��M��Ҷ�z�s�*a���S�n_�G:�/��/���k+��C�PTf��˶���޸8�0k���^H�я~��y.�]=V;�p _T���bݴ<�J� |	{z^x4��ͻxĔt\����㗅��\#`u��m%����a皊�:[L0Q�F�Lq�Zs��b��և�#(F]�,�FVd�A������i�7,�� NW�����u�v�[�1K)T��g�i��|�H�c��t��[*S�z�JRKX�����GN�vmnl�X̵�9��z'�'%�9�H�s%��(��AKqę��U��t�����)%����g���:��3��{���9��Pk^��rb_Y�vb/�Ԙ��G���]a�X�NC�ۀ��c/m����sfH��X���	8��\������0��L��B^�+c�m〰�^lզ����ˀ,�4`zB�P�B�H@���&}?5>�Q�T�=�ݫ�RE�����"-�B�W��6�{+�-����h��W>YPf��&�jR�z`�SE�+[�dA�]��N��+ȃ��p��V���o��i5�*�����0�[^? ��2d�lY�|1q0��Z�@�M0qS��Z�!��n��� ǄBM�&Z��Pꆥi�=�4$��
�"8W�`�b��h���M���DX�1��]�Y;��ދ�3�F4K��_b�<�D��#H[��*��.W;�n�ﰈ��	�Nk;R�}�U� �ԁ��A� ��
�Y��WD��q�#3Cr����V�A�v��&J�&s	6��îq=��C�tI�;c�qvKdo�D�-�kK�eFP��\����$���8�d���yu��_��gv6�L�*:茉4�CL&ؗ��T�%�n�L���s�&zU�ۊ�+����@��1�_�`O�K���7�O*U<��ɤ�e9��蟫��-KE���~�������4v�M S�4Z����� �1 �M"(#���=���3���>D�W���ҧe˔�~���^J��/�B�vS�*v86K���F��D��yɆ��P1�)͝˅]�����$�iSz�k�e/��RRas�4���饡�[%ܕ���͊(��ޚmp��c��5M�J��ma^_�
!y)�A1ZZչ(P�34/g��&yS�B�QRNIf�d%k/e4��J��lN֙騚���d�:M��kk	#v"yAm��o\i�Q�?����D;�,$�3_@m����$	�ˁ�ěڔN��d��P�#��]n�+��� T��F�7��&q����5�l{�ӨO�9I%�oX�����WM�)�*T;[0��BNCH���R�3���+�̜=}#��p|đ�W��H��6������o%�2���;=Ĳ.�>q~Y}M!f�^� ��n�����/�KO��m����%��F�θ`�=r����P�m�5����%?a�[��T�na����.ʧg�����7r�;��C4�CqP����=˩a�gV2�ɂ��!�*��A��\/��� �z�|pD� �.Dv��4�)n�����D�^��}~��I�ɢ���V�%�1�ۭLH�?���fOc��4�� g��<�ʂ%_j}�NrW����L)E���:�I���I�"� ����0M�ǿ;8#�j��J3����݈�1\�Dӌ��^+�ϲ��YHۉ��}6����"O�<�3�;�_���KցZ������������`ʲ�D�U0ys�ǐ4}��_4�ٖ�+X5���" B�j4zi�YP�Ӥo��=4y��RT�2��Y��:2�Q��5ß׆��U���NV�`���||�'Υ��ٵ��|>N�!$���iJ���-��V�J���T&l-e@�Tcf�ٿ2Ƞ/���Z�-ĺ�U=ѯ��^ǔz�����c�>�O%�����<�F����ىn�C"!Y[���@�L�$��o�����묀TK���	|��"��p�'R�_�5�P�L���1�V .96���"�+�)uo<$��+  &���%�k�M
�k���{�8b>�@��(�<!X�z��qNA�@��l8H�sJ�G�IO�udS9��pULd	�x��q�g\�����P�6��q�L�6�tʷ����'%�;��@-D�|�\@}����	�T�*d�r,���:���� mx�k��NLH�^�~�������`������T�n�|W�V��i�a(]��̼���æ(7��vTT�C���vZ�S��G7��* �(�"3�x%�*��&���Nlr/���qܐ9�L�~��* %��]%��휮P-�p���:'�^��0 wGNc��+Ŷ	ͦ7E��e*�a�V��_֎��ݵ�N���z�l�ix��D�5���}(�3��EV?q3d:�Ru�XBn�����Q�e1��$A��7(x%�S�@������O@׶����V��&/P�� ��k�8�z8���mB�o���ݻ����Q��@c=_=�㏗ �O�Cw<K�;�*XC�8���2�NcK���jo��kD�J���J���_�e5/mW� ��B�*,�<���Jr�;���NS:]�\����[���u�6!,�{���Ɖ��D����4b��P'�"��c��J{�!2���&\�Y�ϖon7И"�Rrg;��,����@@�j�0��c�dQ�^��gD��}y:,s9BO?	�ׂ�yw�Hx�jb����I��p��T�N܏��Lc�#����;}�/P�4q}�'d�Cii�ؒ�<���3�<s�A�l����o��Q��#�絜�Qܒfg�^�($��\��m��zL�P��m}�3'x �c��8��L����T/�kc��oz��ha�5 �d5��T�{:�������ou���Df�>4�Q51���I$Ὴ+��+��q>Lkڛ����=;]�L�i��Tm�/�1{@�����ʖS�%tt���"�~s���ŨuQJ�p�cQ�"-�ve'��O��z` ��J���p'�>�7��P�� �i��Г��	��������3��;[�
O.M���u�����H�����%��6��Y�((`��Ooő��dE�ԍ��#~o1g�`wD�0o�B��r���4�r���{Y@>���,B�%�D˦Ë���VW0Z� ��U���
�_YN�Bd��:XK��$���.��ü����:'��g\���C��ۋA{�;�{�.P6��w�'l�Q޳����ݝ>�׋����#z��K�e�0�:L�UA)΋5,N��S�sE�Sg�ic2�'0)���;xuN�n� �4A���8Xzn���ka�����ѻ�R&.rO�X�i#z�ğͽu��B$��S���s;>`����g�X��ݐ�)�u�ݤ���/�[�j2s�>�X�	�Ҕ9�d�~bH�9��}Ѧ19.x
��:役X�D���.v����LA`�L�2@?Z���3�C�+C
���3;�~W�N*I�L-��;� Nru�C�&��;�{f��*�8�~�T�x�ҦW��B�/NG|�\:y��DwOY2L" �ro��Z��?��#����{��,j_�4zJ���͟e�؟�f��,�4B�SS�\]���Y+�{��(|����u��P�E���BM4"�� �"F�;���\=[p�z�+ao%LGQ4�^�$��R��r� W����S+�/z[E5�.%p�?SG�R�?�7cPU"/n�n�=>����;jȅ}%8�ڢ�R)��@����ғS���>��e���-b�����������x�Yw���y��5U�����G�t��J�KW���	���m�mwܨ'�[�ph9Vz��&�,Q��:�2�%P4k1۵MQ/�P$�B��`YھރR���R�<�+6����I�Ũ�f��F4�sn{�L���5ڽ�p(��l%��
*}	��f����;0>��I�ע�)`���x����ħ��lǴ��-g顾`�n��D6�Q���&�Q}�ȋh2��۽M	�,U<�MkWf���}<�.KT!�N�����I���A
[cs�m}yʝ��4���9�r����a��hL)}�u��cf�
[��0	����b~��娕u�7\�$�:w�v��}(�ʃ��t
�.�9)�g�U���>�>��J�>��5T<՜�R���� v�rP�P!8���c����]�Ëh����b��k����`4�F�e�Wc�W��s��,�11�w��ъ�K����P��Y��^Z�2Y�%��y���}�V�mY���=�����dY�a�~۪1�Ȟ)��K��
������Ҙ��P��Q�u��|�T��c	IR��;��;C��5��k�u��;��}�E� '-�J�Ͳ�(��qR�1�h��3G8�Ұ�kH��8�X6�Y;[ZKł?26�����1����9�俓a!�v�U�����4y#�������M�+����Y?��ֱvo��V�8d,�	���x�Q�d"a1��r;�|i0~��� $�6'm�iE� &��K8��Ɋ��f$EPTnHtl�s=F<R�©G�����t�ʖ����'"h�~���!#��s����X��C1�F�&A��#�Z�+I1F�ɏ�,��Ņ|��p����� B���X�&:��ҞV��/�z�DK]�jj��wv�t�$yy� ���W�����H�	��؃Ƕ��a�]E�����)Մ�!��1��m0��掁l�Q�B}��9�y�P~��ܲSΟ ���s_�
�u	�z��&���S�E*o����v����Ƃ�Q�Q�A�C��e��"�>6kB�|���.�k���(��@�{�$��� AXe��&r}�맍G�m���F��b9���7��A� ��P��,��G.:�e���&�w�Uؚ`�Ű� �0)q���0���G2��#�YD��<~F�h�J���,3M�&��g����� �eʺ��O��b������^~�*)��I8����]�<�'�'����">�MM��D.��IEq�����˺t�-��QW��/Q�ٿF�M�q���l�l��{*X�[�,2 '�/�S^ӥ�M���n��9)�3؝+%�4]����p1 ������J�u�g��W��b�^~��4�~�����69�"<���M���еY�$��{�皳ڬѕ�K<����Z���������q�����2Dd��\�g_�B�[��nX��))K3�R���Y��J��y�Ұ�����P=�WGm3��]��~��jDTp��"3Fd=�8�	���̒<�a�����r�8���KW��E2�{g��D<6f;ᬝ��W?�[�W:8R��:��%-Z�T,CC�3ľ0P���,����h-�r���.0�_���3�k;X(�IC��N5����4(���~�'�(UM�)̟���0r�*��b߁jA�`�9"���I���2��N���;���E]��^�z[�n�����t�����7�%x[�z팩Q��旨�_צ��=�?�8Z8��:T�롬����	2�,���V�Σ��JN��iT�sm����݇����+	��Vt��n	�[$��.���C��!����b��f
%e���f�'�)W@v �0��FN�A�V���xV�G/8��L�����YE�z2Z�ru�*4"'�{_gD	�D� ����İ�Т��~��.��^Gyv��@�������S��C�T�}L]����VT�P>Nj'�H�`��扅�L��F�ψB�O�ȊʜIt^"�z�o!"E��M�(�b��B�ߨ���P[�D;-��^s��ր1��<a�b#U�u�}S)!����P�q6ª(��4'P��	oXC$]��t�5���{�>5C����n>c�����R>�  �"s�V}4.���0��J���H���uHZ���(��i�5%��b'���)��/5���ZT�%lT��[�� �����̕CF�T)�W������,������Τ��P��Q�7A�[�t��M"��ʲ�߇/ ��*ft�޺�4�v���:�e
Nrv�~'��UO^?�j#�m�i�g+pH2	O�(����(m�8��Y)>�����y�Q[ݎ�|��8w`yaI�\}�n73�=���+��5\�[���rp|�-�0�!@��?�����t� s:ó���,%�Cԝ�xWP� �_�`�(�f�����lq)�|D����U�%���@8�Z��v������l��G����!@E�n3�1�WQ����sI9!d�U���sR�2K��_�v�[3h���+�Hp��Ido�ݚp���de��ˮ3& ��!￦U+(	������=�6��D����JK���j�q,h���ϑ@"yA��E�IgK��;����~���k�Ð������#HoC�DmB�!ކG��ԗUD�ɘ�x8�D��A ��J��T	�~e�ڃ0�.iXB�bb���X�@�p��5�+}7xӴ�0�s����"pY:�A,�%��6'�H�5:�Cb�<	���	a�[�� ����rb"�p��5���"-�  �2(�g�,�d��B�D��.hD�Y�f�� ~�b;�;�Z�?�_�P �%�w!ƿ$���)���9?��t�'��O�c�����^��REV�F2��F1U@�����I�?�l���=��HW��"�Q��6%(�N���X����}~u
MnE@�7�z�/�n}.Db}p-�_i�0�*��/�k�x̢ ������c�%��Eܥ&�	���T���,#��}�E8�����(G��6�	�P�n���m�T�B� ,�6A��u�ʒ���A�+�Ӡ���l��[l���w?�\� �8b���Ba/��>8nͼ��!s|CNN$�G,�(�k5����F��Dgq��g?s�j6�I&�d���(���sC��2�
���Y?�3�H��s������`��ҳ2�:2b��R��^��u��y�o�rR���fd�T���x$wj�تU�6���r���s��p̈����7.o����,S��4��Acd�
������IPY�}i�ר	�f��ω������Μ|���� fi�Y����8X��06�NG�G������[�.�W�#�n��0�l�Oi�B�ٵ��A�D�ܝ����4л_K^�q 
���e}Rh��Z;�c��������}��@�dR ���:��P��>Z�`h�x������3�C�-l�ɐ۸Ws�Gl�.�Y�̣�q� 2*�G����e��Ǵn�%��Zd/��A7���0*.��RՐ�>/,�����R�N�N�9%B0"]ΥĄ*�uz;̬�GA�%~�����&y2�9����	��^`cŜ�zG[�c;ϯ�O$=��7����s�������˞;-�Q�pS�a�<�P��\�O0G���[;n=FO�Sq� �;S��!��T|�tl���$��dt�,�9�tH9$Ƿ�����P� ��V��3D��m[$��g"s���X�L���!d�a�|�	(����9a:BX'��Rc����I 55�s҇��$S�0�nG��8�.�AMK��揱tyQs0���$=��0�sC<d����kb���9�'x��U3�k�D�O�9�o����+�՛~���r��M�72�s��g�}s�	�?qR����_��������߀7^ˎ0�n�J��4?�>4�Z��ҫf<���%*q���g�/�?�U��Ս�(>�"��b�j�� �R��N_]�8�ɝ[��ڷ�B�m��4�j�E�����?�.^�>�濁��N,0R�Z�g�.|k���9Cn�r>=;,N�g	 � ,L��*ŭ�h��>Y� ��S��v˫�ՇyC@/����v����vz�H ]�*�3{�w��n1�/f������7'��b�������	�RĠ�'���9�4�m�D�{܎Fe�P5���u3��Cy��XxY�H�K�cu�%�ΐ��_�O�,�%��rK�g�]�g`�ڳ������k���ﵳ͘���QǊv�>��昳�B?�?ނ��|f�|���t��|��2��_�-��~�J;�,����ˁ}`����`9�,�����ڿXN<ґLH^�(�^���'�kq\q�譒z�7N����
/����/��5��(K�j݃匭�/���s!���Z�o���t0�I�G��F�	i�j4�O��(�uo^l���kZ��%>��YeW��cZ�jp��#&Eҿr�&��E���b�������*��P ���]�r����Φ>�����Y��N�m������K�օ�ߺ��˗.Q�Yv��Z�!`|Ü���V�xv��@���
��K��R�i�_+s����ex�z�PL���.��^��xd��Y|_�͡����).�y!�
R�j5)t��պ�c؇�H���z��H�M�7,��+���yl������K~2�H�g�M̇z���P�^'E�S�2Z Ah���6}n��MB-�h1:�_N?C d���%�#���}=��������"
��ቪ�2~]?ӊ>���>�]�b���ϴ��
��_D��9�E��[��ŭ��H7dz�d'��c�-��f\�H#0�%k�G�o�ĵ �W�� ��S5����������l"ʦ8(�l��n������|	Ѓ t[��LL�<p؀��Yfmb���ٞ� ��d�����*�C��k-����֓G���j��2Ʊ%.�ar[#]�����~�9�Ȭ�3�U�#�<d�&�D�Z�����R��������'A��B[KWX(��}�\��Z�e��E�]��e�?/���?#�Hq!�����V�@Z�B���}���< ���>o��v�XAVR	�n�G'C�
�}��<o��L%�団I����rB���K����Vt��0��H\��M[h�>�t;��B�n#�^��^�
4���
��u��ϵ���Cm����J�/º��e����w[��Z���V���qư�>A����	f��&���:#φ��|�6�ޛ����@�=��:��D���}��w|��>;1#�6���Хׅ���(��Ks�)���}���iF�<{�cFB4�z�l��I��$#i���'i�Ag:C/�9��c�b�y*�Z�1��t�Y�O�1<Ҝ�s+�]�����麨���G ����ҭ@|���-c�!���e�N��i�խ�� ���+�m��۷]i�Z���O�ӎ�\�i��s"&��wTu6�|�\��O���z��kM�e@�"�N ��A{�������j0��M���#�Nv:V͛��.��Z�T��k$>����O8�����.@Q�����'$0��E�a�H!'������k�Tش��U���h�2)K1����<�k9�$�+���<NeT�6����K�1�*ɝ%D��ӼhW��wjJ��A��L{!x�jЊ΢��;E/��o�)V	{���;5��/�ZS:B�׽tT׶LUi�˻�ݵ�>$�gjHx����\ �`)����|���A������� �� 
��Q�
��!3� ��r�����8�'97�;�J�ٞ�	.fRo	�M�Lw*lw0�yr�Zx,r��f8�`��P��PB[vf�Kq�i(����?dՑCC����wj�Ѱ�3�,�� h��n�H� W�]rf�'s �	��zK���FbpF���ˡy�T��{~8�Bݜ�n��/�h-�F���\�!A:��;��,3u��Yg�����h1d{F�Bnaݾ���֫<qI�t�H	�B�N��.W���*�E�13��a��4��V`����t ��^����M����3�����T'y�u�H��jG�<�M��q��#K�!oA��av+�67�čX�,��!�2,=�!�9 �ɐ���dt��R���>��o� �	����h���7�5����a����Ch�����u$L�F�x�(��E�U�ۦ.�,�Z�-%�Y��U���7+�L�����q�5|����9n䖨Sy��	����W8,C��f��\,H�L*췋D��:�;����N:�P������}Iz�+φ�}�̘��m�j������N՚N�����@���EOD�����$�T�zx�&gO�?~a�}�:%`���\3��$��ZI\�|�x�� y� f��n�aٍ'���=�����mQЎ>�k��x���ϗ3M��e`Ƶ��:s�.��U0���O�6S�1ʤo��T�]��̑���j�:^��v`�+����MGd'�g\�d��	�E�)��������*�P�6�z�{y8Eq���[�R����#����&Iv	�]1ZK�}gΞH ��a/�����B�E�,U?�|����d]���3i����[���Fú|�46�d+{ܝ��u�θ�nօ��*��8�u�`x^Π`������s��Hv�A�&�`�����:�� ���0�6�EӋEm�/8��w��mf��+h�l�Ȇc�&Q�nR-�2ۿ�\�F��x�w��M
#�i���k�����(��NN.'8w>g���?Z��񎻟����-d��`����W������#X��u��x�˭�� ��-X��Ҙ�x_b�FlL s��ϕ]3wĠ��4��1�
0����G�g\�����t�%��jI�1��6���_e�_Ni��D���Z��7٩KTUVi�Y��`�!<��u�\z��Htr��f��e�7�`��1g��tz��������2��=dk9&�*7�}�x�H�|�H�������b�x�0���ơ��颦����a�	�o�CОC�a&AҒ���){-�bǲ\(�d3c�T�{��^B��D8�`�(l���_J����*���4�������4��ޯu@��0ʚ�7|�\C뿱���=���\E5fcY�l��\�K��e�� <�ʷ�Ф�����J6�F��Q_V3�i-� �ѥ�V��0��w�	cY��J�S�L��������&��C�J*�;-,���¢��O��s��Uۤ�K *��9�2�U�bQ�큤��� ��3�
;��$Jh��b}1��_�3K7�_#�Jǿ���E)3����z��;���x+�F�(kf�A�e?���qh�_r�G�V��
��%�5y������X���r���E�\V; ���t%������!��U#��oh�a_�w
�ǨG����&@���]�4WO��7yr���q= *f����O�<I��D`H�u^�T�/hMN8G�hO�w�O|(!m����٥C0W7��������{�#3��7TcL·��@@�(O���,X:�tn������w/�%N(��é����\�����&�S�c0�u�Y�k��o�{�-�I��2��*(ܹ�,��mi��5>i��M�r��/_��w��WZj '8j�U�9�)׷���Ж������k3��pꩠM��,\�d�SPg�����_�VKvkl��ya���D%70���u�jo隌�����w���Y��O}MY���Q
���<�*�|���r���j0\���?�L��-71_� �c���R@p�?ѭ߹���g8'�'��le\}y	�7"~�9�z�}�A�]g&�o7<+�9�ޓ\��)%�*�^�(�����\:�6��֤.G3m�fP��tjۊ����0�7�6�R؎˨IHtAHx���������z�k�q3[=I.�,�~�c͇Q�c���̀��b��J�E%��/�k���pźQ����>�� �>ʨT�1"k��.Tɾ��40�T�M!RHSٕ@�('�M_w@~:�1_�<��橥��k����->��	�&�5Lf��O"�C�K�x۪2�aʼo`^,ЖC���GT?�QQf}��X�����^i��y$��.�*�ń���h?����LM hi"�.������֭Ї��# �m��|lBE�UGl�i$�bw��!Ɓ>4{]��V�̜�/�	��8c�E�^�b�.d������0~� �!�X�2eP�����$��?8W`�K����mx=wl��n1y��ij�z����������}��#�.�@���A!�?���C�'ć�U+F�5��Mt�N��'t�HjF��%5q�@�[ơj7��mtꝎ������FO��β�u%	��f����������������ӻ�\��� �ƶ��s���rXf�U�w����(���9{&�v��rl�31���2D�`�#���S ��a�LअK��2�q�ׅ�s�� H��V%�|�٨�b�5��G>�E�X�����'~\��L��Ֆ�K�6~�D��=i8U���s�c\;P�h~�C��,1�'�E�P�`����D�8�6�V���~ĀT�:���V
�WF �aƿJL(��I�ܬ����O��fxΑy�Cy��� 'P�>Y�˱%�:U 96�j?����J?��!g!{��L�9�ֈ��0i�Q&��p��#W�pT��u�sk6[�x#d-Q�a�0X蒵�կ�����8y��'�Y!�V	�]��B_�v`lc���)g�s�+V�i��و?;/��r��e,�f�\J���P�<בcy���5��|�3���f�Q.a<
xO�_CElM�#���1($d�d�nngv�>Z�)o^8�g���[�!�E�?Ps��\X�n	����Y�J���&�[q�_�(�߳�g�����Nu�g�p�1��_��O�a٦�ƘX�t{5�c��o8O��� +H/t���{�nRf� ~3��ꬔ���=yj���#J�W(�We�= � ڝ�^U�G)s��<���x�B��F7Z�������/6?Zh���*t�	�`lL=\B��i �!�T$��x;znL���7ň������i̣�Z�^���^f5����"lSq������O�A:���bb��&�8d�����.�����[K�]g$�x溕:`7�C�O����pŧZԩ�SM1׊{w-��,�
[��B�����5�u� F=Y�R�������z�؁��!�n�Π��;`i�9��a��[E~?��B�t�>���`�����eu4�hԗ�(q�֦��N�b�֕Ҁ�w�?�ng��&|53r��:ogN�� r��հa�&�E�իl����P`��1l`��u��_~�����U��!��6m�T��Ff���n,C�c�M�v�Q�J���p���]e<���2ą������	.Qc{���Q�@Q����K�R;7�3��J�H�;�� h�����oW�P�QV���b�&�8a�aL�&@�T�MA|�ӾԢ1��9i����d5��:+����q��?�?��J}8�7��c�n�l����<xV��u��+��CL��n���(H��xdr�j���j��H�k�b��
X��-��P���oS`�'�n����>�Z������N��c�A�%�M��t�E��.��n�fMB�i��V�fJ��+jx1E�>�Q�?�d����n�
��P5�Y��"�ų��:����]G��6K���*B�n��~Y׺���W��C��5*?佋n,�E�x�rVd��M�Z6p�G&���(����L�aR`?رp(P��;V��*�gpȹ�_!|2��x	Yt��h� ��.���k�Sk�Fd�?.�8�墶�,\�Y1�f�o(!H�J��ˣa�O�NIˋ[�i��X�U9�Q1բJN�ćѺ���+�}�s�A��Ӑ����|��8P�5H�e�����w���5��O�0���Us��]���h[�Ŏ���+5z6ۛ��WfG �+��#1V�+��1>M��{�X
��9��-F�8��C�ۙ<���w�U>/���$�K���/,u��C���w��Om��|��1q�l��W��r;�T:���nCYV���R4pm�/��Z5��	R��N=K�9�>�����ȓ|��=�o(���#����R7�C�����n�K��h�ٚ����G��4��yc����L����S�0�w�`�'{�Xm�:wv[6~��#]�M���;b)��@�)3 �/&v�"�<�")�D:Ei>-q�>�=""���f���ˑ6J���Gz��Xo�]�_mzo�[H��2__�zgDҎ�"��$�O�!a`k^�*���@\1D��@b�9�Č"��`�>�q7a�,�An }l�F�u2y7$}=1x7H�#,�ϱ�@x8���ŞU�=��y��> ��b���ۡ���G�c���E�|f��Z!f	M��`�c�W2��2�r��%FJ("� tjt�;t^9�dgIc�B�إH���'d��l�S�P^��ƚ�W��h��il6	���۰��h8+9/XW��/�s�7}A�'�(��%Y����b�;������Adc+����p��4�\S��0�O�g�!�����_�����E�����w�� ���9����x<��i�*�U�sixLu�rQʅр��o��}�K���@��%[�P� � ��pl�&��C�F�U.�`]5�_�	�c0�/
����u�Na�W���`1�It��I�����������"��7��%�f2��69A��>�(���ðY�g�6�K�?����!"Km�A|y�|��G+����4��LE�Z�D��S����8`�4C��Fy9��!"#�B|j�����ђ�����Ec�Q#�}�}�����7y�n^�Aa��.?������ȿ��6-�N��9������&�Q]�����#Z5��5�-�T�6'�������G��+�{�g�bš�ޟ�D�����`���Ě�JQ��e�8!�N��O���!BBb�{9X4���&@�����4�V��7U�܁�F�����h��	�c&lB�I~�����E����{xǋ%b\~T�[V��.�f4��Wrf���2��c���u̓lՀd2�G5��,uc�1���Q�E] 葼E��SXZ2 e�[z�zn���ﻵ����������(������V��Gw�m�C:]M�'�����9�%����Sz޽��n���M��F(Xq���%&�x(�Z3p��-�De�^��1��C�ش��e�z�E��=V�~eß%��Ў���1;���3��8�T�I�B+�T e^���pBU߿�7�xxs��q({ ��,/J�W�a�v�#U8�~�u	;�ZO�l�����,�,?),����k͝:ZX�V���,T�,���scy�b����b�.~���e�1��� |W���hV�S �����y�oV<af�2恥��"��_\�X\�$`�XP�|}�^��mU)B0A��8�L#B�g3sW�NCj��`64����/0�"#I�H��m�o��h�}���N�*��SV��FQ�V}0	 C�����.y��c73����1k��3	�0oG����^�0�:'�IN�<Ȼp=���U�-P�d4#�#:q�{�����tˡ�R�m������zf���Q����@�|S4�Ɋ��80^J�o��0.��{�Ό/�v_g�#?1�W��9̘*S��S#"HT�I��� r����U�^ؒ]�G^���&�¶�U����"��^��Xr@�n���iȋѦ싐��������2g�_л�`RO�b���W��hی�:�Y�i9�xG�ێZ�����' t�UՈ�Vg8�3*I����ZWxT����A�z/�a�*Z^Vg���@��se��Bu�\� Z�
%!Vh��c =�X���o�Jl��{�D9r�v�~ڳ�[IX]���PAv�b�yC��������0 �X-�g�4�L��BuT�� �Cyo]U~ьV_��h�d%�t5n1oG��M�쁙o��x�܅pA����M�$�(��iI��_�r�=�F��N��G���S5��儘���O�eڅ��䁋(�A�3��qt���4�gi��X`u����7��/�aY+��0�nӛ����>�I��Z2*��1���É.O&lU��[�Ɖ��r����#[��8!��A9��y�Ԛ���$}YO)/���2_7���p5	G5�PdV
��Κ�P��Z��.���[9��PFT�n=WO�Κ9�řv$k�O��C��.X6|�"m�;��{czce���Z���2�m���Y��N����}�| �'/r�tO��1q\,s��?T�.��~����z�8z؅Pz����f	��wtY�WNe�	�2�f��O%{q�<#i���z�X�7��NY�`�\��0m空�)?A�dI�	���fYu��Jζ�ZX �� �y>�o��"����|g*�z�j 5Xx^��duO[�M��湋Y~�Ԙ1�fQ-S�O�T��������G�૓&�c7Bki;6��@����51ʝu�������)~qP/2���rs��@ ����ܦ6��2ΰ�!����$4ۄ��m,�"��V�lE�w��OFz�m`�v�QnhWΨ�ղ��Cs�X!E��t��13�ڻ:��yQ����w�X�v�F:A�	ՙOD�u .�"����@갾�`&ca-��.��|�_]u�TXe��0S�*:�>p���Bڥ���4�EB��Й�4�'#&�U;hb~b�q�Q �k,�x���k��&�KY�s7'�in�ـ�&EL�Kf8������Y(�����ȼ�u�E��/5�U�=pR�4h���!�7�$`[F�9�;�s�:?.�9�!5�n�F�w=W����E
j������^����'�p�Й�>P�Ѷ�<y!�����Ϙ��b������P��é�N�q^8�vt6�x���TҼ���Iw�۩.�����֓�ZN�8>��<�)�a�u���Gh��Ú���zU}1ں����TM�e��݈�N�g���E�����J�~@pP�5m���T�־��m�^lߔ�Nͯk����� 0q��N�S!\��xc�yʌȎL@ʻ���� �/":�2�ItHg���1٧�u�B��3��'Йj��9�J�Cʘ���Հ&���'�Q�j�*v|\�p���n<��_N���D�Cy�2�2�k��W�t͝KWLW�2�[���$I�9�d��T�x�U�EE����4���A.C4���%��"��� G�i�_Q,47Y$W�!���{�ē��z1�ն��y��Sx;c�~��;\�����/�&Nq���c��,�?na�����l��{�.�l���޲A`���%YG�;��H��陓@�p��(&�bt�З���͍/��}#�x*��F	w�(�=74J��{D�)�X�9y|����
���_��om_>r��2��q�Y<||���,V�����)�l?�'*��u]�J�&���0�i{+���R�[T�K��/�"%ؠ=�Ϻ�PL�p��w�_�/\���Gw�ވ=�<�Ύ��u���s�<�_!���6q�'Td��d!5����wԽ�Z0	��x?̆�D5�ߧ�YK+�TK�˭ y�0wO��7���t�����&��u��w;&>��g� ��u�׼��	}n%�PH*x�	��E)|.�����c��{�����^ ��m�b�!H�uS2�*QОWKl�����9����8�05���A�/��,B��*? �Ё�����n<yə�K�����d4�u[�/�?��B�#%���3�����9�GҰ�#{S�tC0��ߺbKY�0�2���'Si��X6�t�(M=]�3�4T�~������?Kbկ�ZUǑ�R��<��5�k��1��Q���8f�@Y��;;�.�����ݬGqƌZ�r>a6�oY����j'9����G�a���Ɏ�?4G�۩�@���$�n��Ӿ���G:���YNuuć�
xO�p�f.y� z:Q���e��c�q+���ҟ��1�?���C}�} 
>��O���Q�#�ZGKƜ��釚=E��a�|�7�(4n&@!���C���,�[�8;�5P���zT�b]�[�i�Ȣ���>*�f8�K���WM�O%�ǱAP�Y��U��8��p��"~�����jA�7]Lt���,�!��v�N��	��U6$3��7������$3��v��;�a����N��FW�UP*�?F���Ϣg�e@��';������q��\�&z�*G�Q��#t�M����������\k )�g�%)%.2�"a�xY�ý�)�a���%�-l�}4�f�=�۳#�^Wݕ �I�D�A�9�GaU�Hȧs{�_����Tv��������ڐ>�6pl�s���h�$�f��KB|$�4�ȍo����@�C�	Cm-���I*,�5�)��	tR�=Hj�g�:���o%��L��YE���Buvu��	�X�D�;�-�m�>���ѬՁ�y�@�8g'{��	��Qx&�{B��(	� >�0&�����7e��q+H��r4W��4�Fs�.?��	TY���9�56If�AK���fS�^I|ظXQ��X��A�;�tS)�dp��?Z�:O�Q7 0��XN�G�@�'������z��	s=���Ǵ+����Dp)��u��RH�i�H�O��R����n���cux%�iS��oa�
�֞ښ5!t��J�=��"�,E�֩}�Xp�����o/|n��ן[��"�7X�h�rƌ/��u/+6�q��M�^����9!Z��a}H~S
]�����lnAHjQ�5�|m@���쇖'�6�"�B�������e�@�x���*?$..!f�a�$�c@0��w�э�����i1"k��\#�����'^�Gb��cJe72��_����閌ÓwALṓt�;rlw�)�L#�!D&�Ȋ�G@�u���	=p�]��YVf��W���(c-��Mz�7m������R���$�@���GאXW
$�v�Å����C�ϫ�|ڽ�ZF���t�!z��9.lV"���9�.�?� ,^ݡ\�f�	���)$!&ߟ_���F��J��j1Y�$�4���ƚ��>�C���i"mx�c�Z!4�%�?i����� ��_"}i� �gh�Uld9�V:�/J�e��u(��ڱ���]
_��(h�[<?��8�f���.,.@qͬ͞9Q���3��fo��V��xؽ�+�򯞌���gG �V�Ɏp���%m,:���.�C 1+��mw��y�����}$��v�ElO�8�r�Lb�Q�`K�:�����]��>w��l5=����~�.;���~1Bl�y�ES� ��+�SWȱ��z�jMr�Ct�=� e��VOsNHh�ûW1~�����F'�pZyh��8T�$Z�7:,��CV0��.#3�Y����?uq��-�ٕ�#�/օ�qF�c���XutywiI�I�y�7!�xe�}����U��_�n�g��Z�*�a N���11a)Y¨HI��� @���̵4<l����1�m(l(۾����.�P��z�a9wƝN�+�{�5)}~��)��NTⳡ������z`��������k��{������"m�#�4��c'��Vs���7���u`�%�g*Q�MӚ���+�%�V���IX�@������U����l?���ot��6�ٱ֬qX���D���^#��NnD#a�Z�j�3knO���\�O�=�|�|�� |9m��;��#k��#�lջ{�l㝜�cB\�\T�QCŗ��m0���߰,*(��)��/u_%���Q��|ޫ� ��,�{�HȠOc��`��3I;�{E��K��Š�����1-�ݦf����f���ĵ�X#Ld��>����F#���O�H!m�A!L��s�k�%�JM7O�%�Bk�^���9-�ЉW>_����3b�'i�s�E1\ ��sH��M^>8'ya�1��{�	l
.~�E�M"n�q�f��B��Ư�d�y��\d3�<7�G3B4lF�,��u����SZ�W>��p�w���nM�oyA1 ��o�SM��a�s֒����@�x����N�W%�PXn�[����L��{��dH�H��A�r���@�g2����^��38=��>��tt��6�?�S���a<_�Ma��e1ڗ�T0�Ji��K���@�.���g
��=F͵�R�G�($���V-Z�O�d9
L��$s�IF8{r�ĲR5+��EM+�.��ol�)N��6hg���ץK�4�T{>Џ4	����y��O?�w|��%� y��i�I���<Y$+\슴6���Й�����ɂ�ߖ��֡�o��v��Q5��'�%I��oL^0Yɲ,�P�%��p�C��d�]x��x�Pn��x����v
�r t���cbj!Μ���V��c��_�X��V��(�0�q�Ɩ�:k�zN�U��R�:8�x�6#����bQ#7X��� �q�F����l�	�xxl;5�K�E��� ;��\8��<�!aR��'`�U2c75�fgAH�bC_"��1�m"]c��$?P9R�IЃ_m۴���'�$������_���~�ѕaۄ|����ղl@��V��I�����ϳX勈�ܨeUw���[}7��1�SU�gz�}H��=V������Jӷ��e��ᙱ��HV��,���.��I�S��"W��^�T�fb)z�GH�˚�#
�+6;\~�k�YL���T,	�O���,W۹ɦ�|��`	A�#�E=U��0�4���h�<�K(
j�	j��6ZI� �U9�2g��=׎�7�ϋ�f�M�Kȭ%���"��L���D�5d���f0�����
����hw[K�*.�<�uyR9�	���/F;\�$���a�:ǈ��o�}�ƯclmI��G#�sR�09��v^$�{Q�ˍW �ݬ�]�f �DaOK$p
��	:?Z��Jf�&VX�>=�B��9���>)��HH(��i*n媯��_ ���"γn����1ż^��K��7���Uѩ�.\(ey� �ZKӸ^���kA@~j� ���ǭ�����ݒ�j!��ӭ�����*J���WǤ�������H)�tW�"�]=��F�|���������U����Z��d���'·]���Q��}���(�ӌJ<�[U
Umj�}�ۏd1[�@��C�Y��T�W�yO��4���oS���
��]]hs4j\^�t8�d)��W��RK�+8��Ӗ!=�-էg�6��q�Mwk��<�J��+�b���2zf�J��A�Kc�mO\x&��K����h��rn��_t�iJ��(�2�SimW��8g$�BQ��`P<�-2IU�p�d}Ӣ[ǝ��Nt�9b�����b�*����L�[T3�g�3�t+�H�TS�d�Ե��7�~Fv�y���gK��ѵR�5�u+4������ҰW�B���j��D� 8b�r�@��Sc�T�e7^���p�|���KS����eM����Vm�7
s��MR'�����+���y9�T�cƫ<r�3�2(��r�!F�}F6�Θ��P-�۠o��D�+���J���b=�����-#�2}�{��W.�g������u�7��D$!u�a]��5l��2뭮T�V`��w 2���x�x3�`ӆ���>��6̢��щ�1��<�Q)W�������`2�\ֹp12R�(���CN��9�7Z��Z���4 >�m�'4P���z�Dmo��O��
^�����$>�FyCD�@����Ų�s�9c_k]�lT6S�����_���@mMX��C<���T�Bxlբ�~,����9�錷fޱ�ꗵ�v�GVbvx݌x��E]T�	4���;n�����j��@�8eJm�[C�؞xߋ!~8��}t�f��ɚ�ʶ@��dX뉣`����V,�#J����|�xO���
�[F��oɭ��J�6�����>�!�4P)eޡ�un-����'��\�)�� � F�A�)�ϩ=�ҌZ�#p�2��z��G����U'a��βҋI��X����べ֬!��e7�z��>�������ف�������cp������a��`�\���5>5�Y����]�*�-d [<� �=��8r,B��L:����r$�a��Or9M�[��/c��ܳ���苤�i�D9���iA:8��Y���7QQ������T�i
ԅ���l[�h�pz�p=�~��<�dh�8woV������̖�9���YS������̨y�^%�ZA��kM�/%q�g��r��ΠtO]�)���������'9�7�:���q�_�ȌT�
���tt�	EI@���Z�'�$��G	]��c�u1�=��*z�vQ"輊�ԮǛ��"�Őy&`��*�r��؈~�w2H%��b�JGU�}��~](�Ets]��<�o70�)�>�?�j��� �*U��{�\�I��5��7�Kߨm�V����\���;�q̱��������0�4s�R?���v���!dz=Ě�|LO��YWS<p*�Ɂ��:��X8r	ǆ4��s�Λ����a\�u��|✅-f/�_?w�}���0L���=3��҆c�t:t���3���%CB,�2g��|o��j����ow�3ӏ@�bH`u�퐈��
��lY����F��=�G����+L�5�o	DE�T�ݰ��������>���͝n6��y�ꌐ,Q��V*�$��n���9�yrC޿�<����s'�p	��ᩋI ��2��`7B�^�5��{!$��%��mKV�`Vtg�(������I�52� !I3"��O�*laL���x����Nr��Z�u�PG�"���_�>��/'(��IL����.�;QQρ����y�҂��E%���W�Â,���������sajO�۝m�n̜��uA�8�����qkN�P�o�@J��Q��B x
�K95��߷�����^^	�!�p~Ԉ	p�� qGވ�����ͷ��d��tF�;5$�$�p�ci��r������,�2\�� ��*�\������pŚn��"��l�҆���
%ێ4�$5�GӗJo�a7�'s�h�5E6���B��/�U#.�F�w����ɢ��dH���>l��]�����1j� l���P8��İ4��i��P|�o����I+��yl����pG+r��y���l=�|�j7铟[�	6���4ep�q��Er(����� 6�W��-�w�(��Nu�0l��'�c�uq�a��l����bbJ�@�=�_�	hq#��0�%�e?�H�^�]M�/��k8��~��}�W/u,�"t���&�*�ɼ��)� h�����Sy��4�����TLH '��;g��2�⋣��@��K� FJ�3���h&0��_)l����P�$Ӭ���������aR�@�p2؏:4�I���4���\�k;�!M0pFS�>�nu�녪���L:��kG����6��rp_�8��e"� �sdpw����t�Wl�6%�(�Wp��L�|�]��;G��	1(��w#M�qe�}� �.�8��Nq���TD�~��M#���%�!�nVɫzI"�U@��#@lX����)6�.�Y&˕������p�����T�Y`���hC&Ӑ��������6�� �r ���,Qʶ�+�)td�L�m�m,E`XB('<��E�w[j"�����"Y�q�|�Ό�n�<u���T��ԡ�����b�a���QM�����/5�\�k0羣��^�:��Q���|
D��})�NK�B��꽙iu=��Rǯ��Ց9Y�s\�
�K��.�5�xd�q��&�脾��n�yk�\c�9AC*6�n$�w�HE3VV��M��1�t���y��Q��]$��+�Y�=Ҿ�u���/�~�F�{��v����p�3v{n��O�f&��B�7�{p�+���/e��f ?&v�$$%*�:�2�nh�85���0h������q�ɛ����Ku�h�b&2�1��>�G��:(>�Z&�`Z;㻸�Q/�7��_x�u\�Q�P�{�3$\���!K����\�#O)�RS��e�jW�d�<Nn$7�����9��f��޼������yΥ�;p�o.���xm����B(�m�C2��E$p�/p�u%��sDˀJ��9��W�/����-k{u�#��L�B}�N�e�T��~.j(C#G�6S��w�,��T��;QṗC�y�n�rK8^b���յ�˟_�ݵv�y��`�yb�ѐ�]G�֔HME�6Z T�U|T���JP���4a4{k��%V8��(��9�҂�<����
<���� 9Z� 7qS���*�K7Q�%��Aw�;9Q�����o�6d�LZRy��.��ڻ���b0V�Yĥ��!$�"'�ꝯ�!�4G.��hg��_I���%yߵ�aYWx�Q}-e��KQ8�HׯpM��0�B�mh����j�����n�b��oJ���,/͋���h�y=5���嘥nҨw'����cm�3`\�i���U�D�m�ҁ�ՕZ�E��*wS�.��A@�]hևiP��=���]�䮽l��~�ܭb`s*%>�V�h�؈!X��y�@���c Kv4�&E�:4<B����s��'���˰���r9fU�[�s"6�4�	R�5�|�k��1������'�ƥ��ҷ�w\<n�&W��,Rox!��Λ�����y�|�G�cIWc1�׷�X�bz����OG���!�h3��dw���*G�����>,�x�Jw��a"��S���`;��줟�qI��3lL�U�������24��֝�<��E�*ƒ�@L���\7���B�ژܟ�8m�K�ü3J<T���K0����kR�t�3l�)7+�9�$��Á��8�VFmU���(/�Tx��_,+t�*/ՌP��S>�ۑs��u�.Tp���
���ÄV�9�)::�l9y�RݴG�	���v`��Q���RŘ1%����rA��P�Q��)�K1�*W��۽�?�LպoȎ���u�WS�K��閔����!��Z<m2��ź ����`�JSʼn��"����'�n��0��&s���.�o(T�I��*|r���X�8�y�%�Q
0��������T0�^��*%%��CN(]Iwk��=`އ()aix8ޯ�y�R�܀�n|�^��7L�i�~����L�����
�'��B�B��Қ�r���|LE�d�'js���䋾�pv���C�/�
Bj��Q�C�y넆*0���BE"�ˮ+�%�nW��p�7���B��pgt���Ւ�Tדs���R�j"�_=��$k4��?<q���}r��W�pCQ��ÒtK�B@�H�3�9e��L�-{������XC@��"�e�;.�֚��=W`3�r=;��.o䊓7�Nfp*�������Z�TӸ��ȍDL%VN��CP&�X��K��\��_�$R� _�E�w����+�Z����Vk�e��	��x��B��Z�%���@�/scβ6;�ZK�k��n�D�u����iH�Ko�}��oed��)*�x~W���'�A�Nlp�-�V~����G�5�h�`�p?��k�7t�%�@���T�Sq���	f���
gg�P����{�d�|���2�K������4��m����JŜ)Y�g�`�"e�r1Љ[�)t�{�IL���h�(p��U;�Ձ��X�*�o��m+����ӪP9������??�y�/��B�jPN�*
�{�d����>)��g��p��X;��Qpmf��ު�D�[�e
J�k8>P@lm'��&�?�{��Py��7��z�+"y�|���E�R�J���s����=g'l\�u؊�v��:� 6/��OZ���a�����&�Յ����U:��A��.��#�
� ��h��v�'ʉ��7��x�л�tp��a�SˏsvǛ �u����FF�t��t�OsǛ�=8xv�9Ѝ��:�b���ѣ��Y3��jSv@䱓��(�L��
���hb��i%�B�r��na�>e��J��}>c-��T���e
�&�?�Q[����ی��݆�^L���l�/Sg�_�B���Rf:J�U���'O	FM��b�N4�B��Qv-&@�|3,���<�k�2�+�V�����AP��?�l��A.�0��+��?�V!��y���2<B�_�Sjn�ɟ>=f����TݯZ?��^��Utb���)��컰�g%�zMD�P�.G�,����So��sW�؄6��]�h�Dq�ʱ'�>�"HG�������`?�X��|b[ƭ�UO,���H)���Z��A�5�!�}����-T3��q&_��p=���daP�Qۧ7�!I���jU�ࢀ�)��j�� Nw%w�p��h�!cI+E����(�_�l5�%�5���5DQ�M����}�TvMy1�Ώ�p
j���q�����g���,�H������IX�HS�ՙ�a�#��W4X/����6��w��ml����] �Np&�1��m�]����*��T���CnZ>���c��m���v�c����\�c�d2��	� U�sM�W���4-��-�D�x���:|z���PJ��d� 9}�j���;G��R��f\"t���՞��$u%"|i��v�2#��� m�PU�|�n�{�̏���c�������Γx>B�ޝ?f����k)�~����$�cWl� 䓎�U�nRW���U*^M^�0E�-��B�:��L�w�6�B�	��?�|d ��x��G��3���W�Y���v�KtQ�~r���)U���/��N��_Ea�ƥvv.��m>փ����^�*���X��Y9M.z4�S��y͞rbj`|f����~��uԴ������x1"�g�i���M��B�� :�+F�bJ@�k>Q��������8���\ߦ����E����QL2�(ќ[�9��hb|5k^x��&x�g�C&!l�<@�@�-�����V���_�6�+�=�)9`r���w�P��t�[=? �Τɻ�����Q�$�X���.f��;�=���Rѿ�eQ�7�-��"Gi|i��nx{�[�jO
��LuMi[�+��^�Ur_8�Hex��r�/JQ?��FJ��*ٸ&��ER:��-�[6qDtF�LN�(`��\���1��J[��G_�	���� O���*��᰷�w��9m5�B�\ӧ15��]�����EeT-O�G����j5B���S�b��(�.%5
����@��L��`�'���0a�Mp0��~W�wշN��E�@�W��lC�m+s"�먿�}��°���+��@��	vs�v2j����L���)
���w���B�����E;ZNMWWB��'�X�a"P���� �ɟ��KA})k���-�0���{�a���7�m�3�Ž�� �u������r松T�9/?��e���܈��0�n�6�W;A����/����ga���kB���J���@�L���{K��Q;͢/�IKG,*b�so��Nk>.	��� �c[EI�y�;���s�=�c�+xe��#L0��\/���_%�[��Q�|e-u鿥�E3�����_��E��Q���}�X[�'	T#���>�,ٚy����_�!6.��_��s�Wc��N�w��Ѡ����8�r���������f� ۔���lȑP.�m���s�4�������s���(hd��~�����F�`N���[����4>��7��ħ�7[�e���i����G��*�e\'��q�+��o�������g
�l%�KcȰ��I.V�cLY�ȎlҤ 	��^o�Β�=�s��tɪ��36&������.�q�������ȸ���F�-��0���u{Mlֵ���a���-14���3+(x����3��*�
��d�������W�g�Y�	�{]�����V�K���(^�����O��g���0�M�YĐ�@�D�EM ����5�X�A���p���n�(5���'Y�Xh~|R�V��odG-�p��*�z��i�۴��M{	�c�aÏ�S�L@/���}��+�,���*LS������CV)	��D��i���TӖ3Nr��Z֖9L=b�r߆U�&	V±�c8
�u��������j�\T=���>����Ù����LF���+���z��;�o��L�3!��3�Ƿ�Ч�C���1]�C�z�3 ���Q�2(&���.S�ЌR�SZ��Pu��B辎`Za�A�uh��5NO�^%�_������m��N������5K�M_�Bidf�f���N����U�e1Z�x�p���;j���C��gkn�GT@���H0�}6!�W�?H�4r3��σ#g�������ΉBM@����G`�m���'�����T��	�hxR��!��B.�N|B�Ő:�J�u(cɎ}	n6�i�m�7��!��X,<��$FH�c��/��9�oD� �?:��"R �Nt��$�R�^�H�c�g���Ƒ���,���˵�`u�b,��Ƿ6���Jե��V��7KY[UF);�A�L��D���}~<7�5n��Ů�O�K��w���
!?�xj�Jw�f�Ѵ�mQ��p6�q�j{^w�����!�jMZh���F���[��m�+w��አƏ^�h�I�%����}�
"��40��W�����=9��o��1]�LΜ|�Jo#�e@���*�Q��j�9�A�ʿ�HO�o���N@�&H�>�i֎nd޿�G�vb���<]�[����U��#6��<�n޵�i�T��G}Z�xX��`�8�*73<�����*6��d��-M�to/�a�H?(O��!��A	��2��i�~�{�4qe���~�.����*G~���7�Y��F�H�*�g�]��8�V�'�֝���N�Q��`��S�A"}�|�Iκ�cK/���V����.�_�h�e҇�=ȗ]��,�~����h�^?dZ�~��>���oq�it-ɺ uݢ]e>�:/#q{�����^�X4�3�#b��^��[�jp��?��pJ�/���=ҏ.����	�ʸ���6�C�z���	��[l�V&f��T�51M`W�Oẑ���MR�O�þg���8�h��`F�� X��}AsI�'�:���38,�X%-xZ��F��wΕ��nZ��{0�-�H�i뛪���S�r-�<�F��L��%_&�8?�����$PiMg<�ܿ����>Tl�_��@���k{	_��H�<���>�9���1�K�e���W�<zG�x�v�$�HQ�n�륍g��>�������@��ek��x�:�h��"��M�J[���l� �w{��<��Mu��+�.8J�4��`���w~%�?)�lcI�֤`�퓩z��WX��`��i��4w�bG�C�'��?6v��h�K�͟���nL��{z��3+����S6T����O
��(|�X4 8��uG0�@c��((S�]�$qt@�"|�j�))��?�_��8��&�ź��Uc�v�5Epy��Y�f�ӽ3Y
��%��n��;yQ1`V��[Zw+�,��� j{=.�n=������rL�cf��s������an�y:4!{5��=���%���<M�.TL��A��j��ud���K��>J����+�Ft�ΒZ��q����q��H��m�J����˲�6LnO?Em�"!{�D�=%��vK�\h��f۠��яi�mb~�,Vvhȶd��́������K�?����l.%�wPݒ}����%k��9�Tn��@��#u�m'7{�R��/�1C�� ���\���n��?�3�xhHr�fcn��f"���0�dy42���J�7���!̶Z��Ǻ�.ʾ¥t��~S���-ԛ��:7���Ҷ��;1�9Ǭѵ�`N��0���6~d���(8��[�67�=�L�n��(D�T3�����",e�+��#��V��<�3[^ϒ��x8���|��*��CU�n\�.�a�6f� <��.��` �^��/!t�6�.����1�o(��zf1$%9�}��/��:Y&����`Qq��зa�8H�?f�q�)Z�b�?�����SV2��b��ƿ��$y$�-����u��)[ZM���W�4��i��|������rH�S���L����㻒�GU�_�{�C"șw����c��l�;� ȩ�Cgr|�u4�0����8۰O��W�8T����-^��4�@����q&�i$���U��\N��>e�e��RňűKХs �Y &���-ŷx���;7�2�
-���*����#���[��^q��u�T=NpeR4���D$���B`�X$�V-�����ݨ�3��R#�/ix�F�LY4�4��O�e�"Ҧ۬4B����xn�!Tùq2�O�Έ2�R��^�����F[�47���>
OU�f�~,nf3GfU83���a����8y�v`��ct,�9�W�p�c���6;�����hsZ���(*���_~<|��7M�咰{�?\��N�Q�/�%zZ���oY��ւ�cǻ�{��/
��(czv�)�cY)�S�t��[�C��U�bcO�Ѿw��:�f^�3��kD��K�#���~y���������a��B\��ӱ��kH_�1�A��$�ثy?�|�؋�j1O��|���7�	�"�~]�jz�R��Nʄ凹ǣ���O�U{�q5�~X�cv���
S��j�!�).�U5y��ԥ�^�$ct��\��-ʧN/�g\@L6"�l���ve�T)8�����8��`��W��H��<��>��Q�]m�ulB�[F�w��_F��,	��M�$$�Y�B�@ W�v�]�� &��/�T�N����qy}Ja�,��I�A�r�tJ�V3��l�Q}�#��V��*��P F�18��X�(.|Ó�+0���̫����1�����~	��H�-�0�w�-4�&�,�����������`A�y@��w���TV��)��_{>�C�n�~L��d����e�Tx4m�!��B�_r���\-�s�mR��g��r#8��������0٩ǁU�,��V֛���Y�b,x(6Y5�v��Kk��[�󝁜�} ���0\.��X&�o�<o�a��܂M�h���MW&ڜq��Բ2C�"�ܜ��nA��u4��7 ��M=��yx�A�0���Nh�U�9�r#�4[��}���^��(y���@16��<�W�����OF:��Zb��I��=�;�`��4�V�څv�N9t�>tEm����!�D
�3��3��c�(&�2qD��6#�/��2���C��H���)��F�*��ӌ����� ��.eb?׶��[�hr&�|zrU�0��F��Kc�O!ru�9ل;D',��R��u�Ls��s���x��\�U��Ӳ�p)�/�"v�v���!�~��Xߎ!�&��Ak�ɨ&7.���H�}6���M=��k���ӦL����4(�728C��3vA+�_<[#o����iT����E &�AV`/�EU3�Ɏ/�=:\ܽ����{�~����Z��"�R<}�
���%�Y�p˓֛z�Ҽh�����=��z��}�J鎺��S�82���{�{�^��5���E��m=il���Y�,�w�f���HM��y[�ds�X�-u����*""_���Q���K�HF��l��f���4zIl�x5�λ|�w������4(Kh�`�>\� �!�U~o���q��m�����<��av�ǉ���W�Y�A��a+�x@��k��=�bz���[�r���/)`K'�mB'��h{�\3��-!a3#DI�vSI�^ZAL'���^���c��E��V3�LBH�$����'�\t��͇��I9{�6�9�$���,�Si��ATS�8QR�a�1�����y�L"�E���K�;�+�*�r����;��U���M�wނ,3�{� S-g�;N��|c���~�,ͽQ�ә��b,v�G�����z��Go��.^y1�^�X;y���U�Jf�+�B $��~�\�Y~�A��ba���h%X��o�mQ~||^Y�ʈ�xu�-�ڥ��J�:Z/ߊ�wf5k�l�S$�}�*�a�@mEy��XV���})H��Q�&�)����L��h��O��1p�=�8�k��_��éٸP������)��{�6�:Q`53r�9�H��X�����G��!F�����/f
I���z2&SB)ӑf:z�`E��:������-�6yA���6��#:�*٩��*�|���&5RL�{�畼�p��Nd쨄�T�LI5, ~T[�&5^�8&Xݼ��7� �Z��c[OA�Y�)����H]�R:��,�)�_�8�F���)��B��� s�/&s�Ώ\�������=�h́�*$�]����9�Yn���-�࿠�i;�/ �ɉ����\��*|�����[sK�O�t"[�A$��M��^�yv>,����,#��~��[X-�I0��
`�Ss�OA�����x3�O�,|d��44_��C�����NMY�i=�y�Gz�`p>U1��u�z�6���٭�������<d�rInb�H�-bě��v�����7 <H_�)�*:���X���$]���OG``��-=--[��o���\�������<1͆������>�������r2��}�۔�I[��x�5�_�t��7Y����_��Y��O���i��䠅ۓ .A���m��ޫ�_���-�	�WY6�L`K]��f ��C��&��4�?|���H�x:7��\��rY��(�~;��c<%m�+����|N_Q�P�N6�7�q����q��]v����)�{D�Uh3�
�m!��'}�Mg�58L�F̯N��]63�����ɱ��;���딄TKڇ���l�C�����5�aH�T��v�h~f����'������5}˴S�U�Z~��rgw�P��
�h�����|�6E��h�(�GXD��;Ɵ�)��m�)���y�h�k������;U��X�Z�.�B���>ʥĔ��O�JeZU����c#���Z�!���|e��[/V�������h��f��D#��ij v�C��n����T+��?�war��ʠ"-T?����R�]��	22�����1̶�Z!u6��������Y�/��C�R��j��p�R�;0��_�������^�%�P��*��9��3P8`b�%f���!��F�JN?�C�S̅�}s�v��Ou]I�T������4����w57�c�N��v�,ܶ1�:,�j�.Q_ׅ�yS��ĳ���EZ�1����-���
���*~-�"p����0`&)��W̞4����e�D_��k��b�%������k¤�>�ԉ
���R=�B��?1�7�~�w[֌��Y���� ��R���Ps�Qqw#n3#6Wx��Ua(�xlH�e�sS��'ϱ�͔A���Ԅ��$q��v�����%���Ԝ�y:�l�`���n�4�Դ�zf�B��o-S9���Cj$�l��ϷP�{�Ѡ�@��a�����K�&���p�POcs���$� �6Z��� 2��,�J«UYI�'tA�"͗�����l��Qi����?�k9���u֎���WN/|n#N"����3�ٝ��:M�վ%b�a�Y^ȕ<����6��\x2Á������!���T\,��+Qi��@+��l�[���<E(o�4],=#)����\gL Ģ�G(���D�'Hx.��݈�׫V0��C����[�����+�C�3+|w^G��N�Q9��҇~�K8�H3�|�K�K�hCI๛,�l�F#b9���E3ɳ��N�( ���N������w>,T��ĩ���ej+�{��߅z��$Lz3�c��tb�hX���h��ŀ!Z���f�&ƯS��L�};�ҍMf�NBb�dP�#���s���d�7�`���%�]J(.օ�҃8נ�:9�߲�����p�Rq�OSnb��G�F�zp�F?b�߼���?6����MD���*:1cV)yD-/���)��n�tnQXD9&���av���v�H[��'-j���b�9)εRb1�����Ra|�;*��Vچ�\���K?��'9�φ�@2���6���?��N4�bV�Z���3Y�<���r<�3rQ���v퍲�s�M��G9u�@>��h+@�Omz'R^oRe�#���״���2����/��ȸ�s��>�$��M��|��މ�
���B>7�Ԇ�s~���OUeaV�L��+�k�\�eK��Ms�v�yM�`&�-*p���ã��ǄA
�rr���?[��?,����б�{1�������հ�3�4��)�q����Áz���)ǿ;OGO�Bܜ�r��qxsI�Src��_7�76&i0�0���N�iP�����ŅD�#�K���;�I~!��i�5g�c(yvD�� ]�]�b�Q�ɬW��4�i���h̊�w\I���H7���O���Qs֙���uc:9M�������\7��5����F��ʨ��ύL�%��0s��14mޒx��l��v�otËУ޲�g����
�|�J���`���V]���-�А>�u4����wl�vy+,��i����x�I��j�����L�E�K��Cm�֖��RS����\ 編�U��z2��m�	dcOʔt�$O:m�����m�)��<`��mq�i �bBP�{��>uE9҈��R�ק��h0��:�,� �&���cq�Rpk|ќ�N��ѥD̥< ��,���@�a����V.���`B�덄~�%S�+�q����a�N-�4|e6F�RZ�S��_��zְ�:F�&.��x3D����Y[T��Эą��{���nǋQS���Ń48���w�o��\��͂
�{����K`��s������m���yEk1�v]�N�K�p�`�wL���F�Y@@�2&��-a��ZO���B�H�� b%���SI��R!��G��s}<߳D1���E._d	�5c�a����?��~�#���QkYU�AG)��>�����1/P����/)x��-�"��0 ��-@�E�r+���:��(+Ρ�|�ʯ���;����� �K�^��I=�E��,�-D����_��FM&���a�vf�yI��s�d�j7Oi�Cv<�35��Pŗ��J��S�o����d@!�ʓ�� �<O^ۛ�[i��R���(���Y2 B����] �ӣ3U�{� �3��\����F�d�hD�D��-M;��յo�a"�Yh6�����h�8	R9\���B���)�X��h�������>�I�&6�E]o���ج*���s�C4�@,��k�x����]U��W�B���nk���n�L��^���c��-p��n��V�j�3C�� d��s��������X��Q�IU�t�)c ���|4�!�d!,h��m,������ �����/gyo@5���l[^LJ��]ҳN��v���m�\�&�=�4��p>�W�z㙇�����ڔW�eJ2,�����w���p�	�p�f�n붰����A�EG�[����D2u�U�;!�㜅����o5h�#8�4��+cRB�76�����|�C��{��AhS{R�Z7ɗT�� Թd1佹6WQ�O[�{4YQ��' �0�Z�D|?����B�dwt+)��L.�zw�(/[aY2nh�_�1���S_f����s篇97N2ly�ڻ �9<N�}��!��ҷ8y!~;��ֽ	��SӚ�+~��LP�D�T��/G]j�.�"���ӯ��� �<,�2f�x��:�#5z0X�3zq��.EK�����'?�����"�n� !�r��uw*j�.��� %bl��5�}��m68j��O��qt��}�iI��z�����I���&�ԖzeԌa�KKK�ċȳc'��`]R�]�K%˰����B�fL�('m������@y1��Z��,S�&��3ɻ�'�l���݊�R70[:��5�Z��
�	`bK���.>Y�pp7�b����{ܢ����v�6H?]��I�I�B����չ �tDeDػ�Qb�NZ����Ջ��k���`��=T�wT˿k/?��G�8�5�FC�y&C�5@�[E^��ܕ_?h�l�DRT|0����T��s�S ?��-�z���y,�'"�к�>�w�-d�x�H���+ y���~��+���"f���y���Y/�D�-Q�5yI������{�Q�Y{���
_���q]�$g�)�7mӋ�`�ol���Ae���gi#Ob�F@����u)#�M�S�?=7�l�E��f!�gS �zK���
s�z]h='&����'�01\4���F�3���٫�DR@0�U)���^�t���>�u(l���v'�kt7ƛFDG`���ì�h�Վ�^�����s���QW�nV��![�cq\�7��4��
�Ŏ3X��HI�Ѥ�yh!�h��1�e.�Q6���Xu|h7�Ev��ſ�ۑe��~VST���y����s�v�����?�H��Ra��J�S���(.�
�.ثr����R��џ2�h\Kջ��T"� ��(1���d܋���]���;8�*"�����fd���|�����+'KM�����&�_���1�L9 �n ͟V��h���etm:eG��x���J��s��˅�
΢S���6���tSio��t�c�J�!k�!
D��8+��0k�O��('��8
d����Ne��I��^�r"�Y�6j@��N��V4�0,h�Ȫ<�G����"���mR�V�1��DKC��列S�?Wp�wJj�a�B�Ԉ�-_nVĀJz�����=�tR�� ���Nna�֗�/̩�/��P��oc?��Z��9٨�r��ۃ<&{(�q4$,�����R\�+;y3��58�<+9��i�s�H��̲��n˝s�z�W֎kяo�U	��Czy�|�uƺ�id��ju����PR<�l��9g��9�������,�z��3t����c��9(/�<�?��ڨ����	HD"o9�u����u�1M��.i�L��oubb,�~�3�B�P���݈�(A?<{�۔i�m�A7�%%D�Q��z��`�/�n��|/36ޖ%|Q)>E�ZuI��R�W)0��������%炘���^֤�1��|����T~�B{��5� a�����˜b�{�D�(���@����_�t�����r�͛���R+z<�h�fu�I˿�fo/��tЏܟPP$SGP�qLu���=�c$V���s3P�Q?Q�`��y�a��L��k@&�����^��uAj�����}l|*kۆ׬b�WO��V{Cjj�+YRr�Z��0�}��d}>��,XRz���s�����¥T�]�VA �3��ԴA��tA�\��/��c�0j�9���#�v��#ypi���6��!��J��B�Yo�b$��3�:�磻:�����Xk��G$�
w����j��x��!���V�����:dLm����^
�Xq�2��O�f昫;���̼l��J-o��KJ"&�}�V+F6o�C�� �	�m��cL\\����<n �j�f/n����T;%:]�[`��h�j	��1���u���x8�,��&y�e�y}<s�fܴ��d��$��S�~�	_J��XN��^�7^�Q������y�Ŏ7������\�e��'a�n`K]����f�;�Nba)�)�q��/M����U
¿�ENaz^=���z74 ~8e(8��nX��O��{k�8�ď�zb�I���&S���βI]2wYA��I:����I���-�ZV���'���WfW�!���Jr�R�(��O�Ƞkyd�4Sx I��ב��{�� �ݪ��W��eH�H��lp�&�仹���_}X(r�.�עK���X����Ó��t����J�2�'�c�P���ݲ�J3��D�2ٚm�9��L^����E�ix?¿+�������*�A�^��Zcژv�[�9V�/]��C 6i�$&�ZC�������4��c%?��ϵ��{L���ol�K�9�-*����:=X/����K߽��WjP�i�]o42�N��H��rg �P��{���<��o=�è��([5x�=8�i�-[��x�xp '5M��f^��G����4��#Q5����
@t"���:.����Rg������'}�t���(ʳ��_cX�n~��eA�B��~t\y���U;#��\4=��]Uc&�
��캚8#��>k(ȉ==�W�`�|p|F셥�{���^g�a���t̳)V�� �E�)��A�B|7�pH���{����6K=r��\8Ѷ}Sښ�8�*H�,�^��E1s�X�Ge��]'zr|��HM���¶�8k*1��6)�l��S��O	9�K�]�JU�k}R;,��ZA30���v�i��߂U�bi�_O�#�V3t�]A+8��]j�z+�!6�o1���VÝ7X����y�Pz&f��*��(���ֈY+�L;��R-bp��ڡ�@��O���bDA&�y�������1i����	y*��K�f<��(�!두i�M�Q����د�)j�oB�k�$�o�t̚'��Y�eTcz�w:˘m(Q�gӦ�:?c�����ݨ��v$��/g�������F#}�����}�O�q�W��a�5D��T(��0��~6�G���
����wJT$/�χ�jzs��S{�q��Z���e�d�*��~� Wr�3J��C����o5k��)cE�bȐ��t}HTi��ۖ�e<��{R�Je�]��V1��XU�/2$���VOjZt_�d����5/��ɳ��A9EL�
�_�|f7�Ѕ?��F��]�����;B⃤K��e��_������e�i����NK"�ʃ�
����o���,��y�bnPjp���i>k�?�j/"麗��>?�#5��;��O��h�9G�"�tsD�X���jo�@R��ϖ�!G��#Ѩ 1d�
'�	�I��X�j^�����)��p�3�.VQe,�qw�;_�r/��K�e�,���/᙭�/�����a�:�=ɚ���$���X��2D��c�ɉ�� ��$]G��Ei7.�nc�vX�l�:H�%�JJ�}9�C�&#�2��ѡ����d}{��"���xc�Sm4 PxH�A`H�v3�0��b�1�Zߔ4�A�bj{[�sTј���tL39��m�	�7J:�	�L���]�^��
�c�"�,�|,�<��$��Cf���3K9 /�4�TGI��VD"���������]��e�1IkѴg��,!�U���-;���u�|�p���(c�%��O2S����GXY)'�t�H(t�
Wx���C�f̉J�ï�ꯘv1ؼ>xm��z�5�Mw��C�u;0�L�>�7$>���i�0��؞׎�[��.(-e�zFF�ű��ȿ���O��O�pW^�=('�M��k�py�F4B�ay�3H_�����H�{pg| �����������˱Xo���G��^��Ã�r ������z�4<o/f�v�}5��)��� Ĺ.�Nɝ����a� 9��*!��#�l]��.����Ѯ�B6'�iWj�)�\��ػ���8�Tp�����Z�������X����&� ~pڳR���^��\��_R�`��NY����Cg���(��Qӈ`��l�z+fٓ��E��[��v��9*��B>�%�E�����\�BJ�Y4"�ޱ�@�[E���0T̍������7P�N]Ζ�����qU�L�fG,���<�(4�\k����9�����bD�->�"�wlD�4���8��#Z~��ec�R��GX�52�ߘEU��5P�O!`_�r�$�v1z���/f����ǾJ+�5�����r��֍����$��g4�93eL�h��m��F���OO�P���U�PF�ҹ3!��Y�-��`S'�K@�)����/��N{����4��"���a�s���|)������A�حʞ7K���<D����d�<����;�E>�	�${y�?!�G���U�ƚ�ÐQ��X�IB��`��(�tws�}N�a?�)�#bݓ�Iu��Th��sH@�ta��,7%���|*�0�h�Z���<�I��)|.�`3�9�dr��T��ֈ7:ȡ�<"}`Aj.l��.h�t�X�K��aV��]{�D�����u����.���2�Vj%VȽ^R�wY��b8�@)���w���n}uQ���/U��z�l	�_�c�jt�
g���t��H�4�#פk����D�O���c��`�q&���g��X�\��6��@ƶQ���N��b5�v�*�.E�~�����Y��퍔�P��s�H-�>O!�&O��DI/QF��i�|���Zh�^����
�|���7��e'�?=�t薊./��hDv ��[�͵]t����4�c��|O���tzڔ�&�h�h��B4��۹ԪYų��ڂ[��(`�;��ğU�f=��cz��u��p�<�8�'�����d���[�t�f"�p��"�kKТ|yg~-G~��z"��v�co|E�hVM�Eh�V�/3"l��KQ}C�� �WHO�[��B�WK�LHB[H����HWX<�\@��9Tъ���6w^BB4Ӊ��lH��p�5�ɪ��*r��v�ўU��d���S��
�a�'Dp��ɚ>Dco��@��/�U��]�p��U턃\��KKe�YX�`�2�Ν��3?��c]�\�,od�)�2�g�;���a,��y�i\�=R����j�=��!��oZ�#��y�f�����˧�ٟu�R.�j-:��<���@��TT}�F�w��7�+jy56IZ�Ѵ𼀖��;��]��3��=0#c�:m�]�H:���~�� vDC���ج�`��RfƧ�J3��m2��T��s���1�պia3�L�����7�2���������r����5L�� ~���b1Q1��=��!,�8�\*{.i/fڰ-��j�n�
��V�$v�������%�ʓ�N��0����R�	�I�2�5�g
R��aAi�Y}�^<����!��S)�(c,��Ψ�:���D�95ۭ�T���d�T�M�3
g�ܚ2d�x`�(��$F��Ǭ��d�O�h�%9�=�D���
��9D�����q���W��db=�M��"��pƭw_K�3e�������||uL��'�2�����[��?[!M�&ڹ�� �2�:�����Sfa��T`�*���3��~u�c�2�:I��R��HQ1{ �B���FYKz�劓'{���sJ|{�vG_�xF�� ]��r�����g̰�&z�&=O�a�?!m�����W�G��#u�+��(|����:X �� UN ���P�L��f<w�f��-�ov�_ר�P*<U�:�%���Ir���{�#���
�o,_e\�Ha�sU�Z��>5n�|:��K)�m����K=1�I���QL��^��$��	��q���S���$���J�.��>�g��Q�s�h�v�֪"Rg����m���w֪Fۗ�%&������6;�
!~ޏ/b��e�Y_����u�p3��\K�@�4;��<<�!����2�������y�0��:6��;�K���I��p����y�d�ӝ��-�1�� ҃�)o�*o�ՠ�=�;��!�䞕�At�o�":��*��vk!єz�%���&���c�*8Ko��9�
K�Ɗ%�R�
�������:�{���_���j�9�<Frka���~��J���PToK�L-L����a����1_cܱ��A�1���MpP?-l^X�Ȓ�6�?DLƌTAl��,(9�$�1Zx�x��r�� �
+�tF'0#;0�:� h#
C-2�s]IB�Y$�kj.�_d_Xܲ~�S`�(��BU�%��.����ŋcJ��l_�년r��|4z2̘�T󱐀�O���5��X�vs0��g���rӠ궯�O��	��I��P"��$/��968����T O��,Q��F�yșh���NH�	:_)�50Y5�&����`�8�I���K�K�;Y�lZ}"�ݛ���:�>���}@���_�@Θ4��b�#��y���}��P1�He+�2^8�͚�c�K褷����J1��}�x.w��,�\ZTL	�,�4,_zd��;�b��yڥ�YwX�/�s&c�7$��:9�e�Zp#� 8n��	Fc���%��A�z��pM��콖
�w�߈��;�� -��h�������y��|s�=���Yzhm-V@�$!��2��K(�&Fe[�-�&�=�P��>�R����g���n�;$�	>�e�����w���ȶ[�>�����Dcp�Y���a-,Q��="@�2�?���ՠ�XU\|-@ �[�͟�g���L^c4����uMj
�&X�@D~HvW�{�A ���KFOO|�	̟GȎ�3&M���Vh�,����Y��m�t��\pJ��l#�r�KJq8��A'tP�#�̚��.�3���(��p�|��}�k��}R�8d�����?�"G�*b�ze+6��di�DOfV��@<TАj�x���&�m����H��]#(��Bs�τ�Y��it�AE��ʑBu��jd�9I)��j3{SKr����\������ǿ�����_� �&���>���;ß����+�<C��&(
ųK�޽3�j-���?�A�/���m&�|<����W)^*?�M$�����ھ�vcx�߃��{Z�
e�,�
z2�Z�������_�b���]�G�()p7\�/�?X�B�þ��\���ȴ�N��YK[tW����1��>z�^�9���	�r�����J���C�[qe*MrSs]G��%\,u�;�v7��Srİ�Eȼe*IHmB���~�S�Yi�@T��Z1(p(SE���0�2����_��)��#9����hz/�b�����0�ڄE���Y��)2��2���8��e���#7�~��C������Up$�R��Uj9.�De#TH�KsfI��<U���,���*P�k��!(����d6�'���X�-�n;�F���5s���*h|M�e���L��},B7����0F���q )i��H�}��|�zlka�� 	��zU�;�GM۾�D<�
�$9Pj�E�v�E�y����"�P�Q�/���g�i�K�E
-�������]��&���۟�[����3���#��W�I ��-��N΂
 ���c�z�pS8����䰝�5�L=��d;�y�zCN�&l����'g���M��8�.2O��"�mb����RV���v!�:��9�3��H���Ya��fE7
�m���D?f�{�M<^���<ԏj����a�����`�*|���(��rO�_�{���,4���(S�{�^W1�%���́HEyN���3�_�$ޗ�0Į0��b���� i�1���jL�?��v��y���r�q����XES��'���ZM��C�qΉEuy`%�V����]T��,�����Op�Z<9�)�L|��1����k$&�����5ʳ��X<��$�{yJ�r�&��	$�gn^ñϭ9k��Yq�~�T�P�<���0.vU�N�j%�����8:d�7P�d�"���H:,���>H�\��'�i�>�n�1��֝�Nyy�I�ߏ8i�����L
��.{��F�TW�T�*��/�����n�I�7!�@�S3�!���2mw�Qm.��Ɗ��$��S��on&�k��m������
�/a�j��0L��~ w-�����liZ�at��>���GY���ܿ4j�8�Am�_��X�!�L�B#'���E�m���5������&DI���Mu:�����a��ؗ+���b^�Ӳ:NŎ]�"BVtM� �ֺ�1�Tz(��6��:����i����XIk|���A��.�7�̰/C��[:����м�>�0(�%0��饔�e��AWs�*���<8�߻N݈$�T���S��I��[�Ͼ�/Q� ����`���	q)"}�G=�ף��!���������#�<ػ>syC{�`[iN�wW��qG������6��^lݠ�Za�����v��H�%��W�T]L>I���S�գ9�"��aD9ެ7�H1,E��G��5��V��ۭ��\�A�TRjR���y�.Z�G�Κ5	��S�W<��ؐv��.v�P�;��`y��ٗ����,R+\�����U��ƶq�p;�i�FL�
��`��
Zpʵ]�r"��_����+��;wy��k��O�GvwA� �WM pM��+s���j+hYhA�����m���~8���j��	b�a�thCt�2W���
��&h��I�G4�=��a~�s#�l�t�p�2g�a��u�7�
�́�x6��>M�׵yy��@�i��
�i��)V�@�!C/�Ap�*� ˚w��b�9l6���t��ۿ&L�5#��5i�;�.�����ܸv13Kԋe/�SǕ��>���)��JUr;�o��h?J- � ��e�ۀY���4M�ٶ�����hz�}��t���e=�j=p��� �@<"\���i��i`h�@�����(��8�F�~h9k�t����7L�c)�x�!1X6`z�pD��䅴���Al�'�{ċ#"��=���n�؊2�is������Yu�*P	j��)�|�m����_� A�]��)x/� %w�UHm���l}QK>P��Ug_��P���2�:�q���M>Y�AѯRK�Fd������G���j.n�@.�^�?d� �O_����h$g�U`{��۫򊜀��o���g�;"*V�V�[��!+�a	�fǢN�ad�ߑ�וt�m�~��D�%IJ��A���ZyqYafU7=�4R@�vMm.8��m"����U&���_sDY�3(U6`�*5�Ys|��E�� ���0�Ә���Eڎ�떦�/�p�Q�mye5�0MxRS�����J  ��e���U�o����^�*'������Z���O��d��.���RԚI�|��ij���EYoC���iB���Ɠ��d���|�<�(^MT���h�=��O��v,ҿ�r�d���~�(���V[�E4����(��Y�:�;�$�Z�0G��o�&��<zi����K�
�A��VVj�x2�Y��R��3�Wn��Y�� .ݳ�U]�)�m�4���ۃ���i�L�L6jZ�uO%eq� _���Wfg8Vl�7k�ͯI�a�o:}k�'ˑ�6J�wn����줿߹$�SK1��~�֞�����,,���J���wB�ƺ�bZ�0[�$�Ow�q�^��T/>T߽��y��X�[�)�_�÷׵�^hn�
�T�6�$��  y����!I��Nֵ`��z�+R��<xEMbz)��M:R-��%E���W��S��׽1�U~Q��$)_r85t��@�R7�T2�Yg%�O�h�P�:>��0F��K<cۧ�n�F��-�1��e�G���ET��$����j�V��Y��m�����߂�fIc�����i�)k>�����Fb���d�Z*NM'�\� �@�=59g⣞P0\����t������6v��<G������w���
ޘ�t�AfH�8#FA'�D
���g������.�A��cr@���BO�䁃��C����O�8�w`^(��e>}f���X;
�,?[��M��0�p�l�Z��a�?E)�Yn�t�S��}�~�7\�*~����u�CE�z�#�,��7����W�5
�3zc�3�Z���ٝ;UOe��-PT�(�ҥ���X�j{��~�4gY�e��+y��,����9�۩����F�0��<���<bpQ����F����!o��<k��t��N����*1�Cg�Pz�f6C��E�������Yp�iJ%�@R�Q���s$B�SO��gVo��)",�ֳzcB}iq��ye'_Տ�B�U��sᣳ�$B�F��gr0<�{�-��6	���`��5�6/,c:��B;�.0�.Z��Q��kE�%�VH�	[H'�I�6Q`����*��i�_��]�ɕ������ϼź�VI[Q�v�i9̽���md��+�Ty�bF��hp.��z��ǻq�s�}���Ae֟��ͯ���e��E�����K���L��ɜS��Z��>11��l��b�K�n!����u�mCY�^
�sE�^2|�M(0^i_�������[ �߿}�K;��z�1�-H�g�\���{-J�6`XMγ�wL$Q&�'���Y��:�	�[��r�3Lne���U�cW���l��U�U	R*F��i5�
�������P���m�ߕ	*VIɖ�}���"����nZ��)����;�9D���D-����^���R1�������:C/hi7���m`"0K��K�j�����B�ptI.%�t��>���^M�wLʹ�B���Xdfӫ�e�(�?O��=�;�Ȭ/J[�l(V��u)s�w����W��K}�
��ƶ)�+&�8�V���2" tv��Y������Y�o3��[ݲ����,ܮ7����
{@n�w1����SPN(�-:o�ZTu5`6Ȉ)X.�� Vs	+���4q.�=5N�Xpn7ױMd0wCo�JØ����"�u�3ϸ)��G��6��L|n��cN�ڊ �'ы��X���d�L$t���YB9�?<V��ÎS.��΀#�a�����JV\	�x{4��ل#��B߉_��g�j�-G����e&ƨ�3Uj`�k�x&�ݕ�ƿҷ�MO�3e���E�{�o�6���D��`�z�k+r���N���W#rdԑ'�T�D�8n3��l�U
��h^Î� Mj d��V��W�[��*��[ ��F����9�t�Dd�\xTz
�)u!gu3�m�3�ƏX��t�ʃ�BDQv�H�\C�mo�3�@K)�ߊw�����p͐ύ��m�{ϯ�������8����HT?)����2n5�>�KU 0����]PQ+*�_�Os�oZ���k�X&�`�N.���7ȿ��j�~��ٵ�NT#{�Ò��+X�[K��瑱�C�mz��
�Sh�
�JOW����q�N���$0�bV�s��]E~@ICFo7|4*�6l��Lr�vy�GD�uBi"o���T2��O�Gp����3�H�s���Z��<N�A`�*�mF�k/#cބ�e�"3	wpc���S]o��DxB���f
婵�r��э=�%�x�:���@9�F�p�:�kݯ"����kC��{NM����Ҍ�JG�N��l�u^Vz�X����� ��?�����_���1װ�V>b�Ų��і�����Ǯ`���e���i��^�}b������T��.���Bt .!d�D�~?�7����#�9��ݧ�B\�"�Ϸ�{��fYp�|/ٖԝ�Hp D!���.XZ[q~��A2�(R�[�v푚��_`:`d��ю�>j\��u����>!�H�ӓ��t���,����7s�j/N�;A�����<C/)N\Bz�N�S�ϳG1i�M��Yq:y#.M�.�7Ʋ_2=��qD��zW���m_-��ݷ�_Ƕ�I ��DV��"������ӠґwMJ�Y>�,v0�
�+���3�����(�q��YLȚ��$]Q6�:ALj�r&w�@c)�D���C��1��k�y��:�y=� EGK��������'�`��N��~�95�?� ��dxυ�����n4*���[	���]כ�g���	��\Gp���`��{
����,�@*�*������?���dĐu`u�MJ�]�k?/8�!7(J��/���u�Q�p��;�:�Ē9!����G�a�{��._�ߣYW���*�i�b~��3��PS��PՖ���_��,�����J���!���a��a������Y��^>�IV��5ے+��)�X䁵��<�D�5�w��Q�-�;jN��r��<��1���:a�2�f�� �I Z�
)+�-	e�b�h,K�����v�����
�_E;���[/,+�)�c1��0)�Gx�!�H���J�2��I�R��.�l����O٩�R�����f)Z��t�o��	����w�0&��^ķ�!Hw�'F�2�8�$8��t7����MO��C�rdv�~��h)Z��b&S�?y;��c���9�?n������ë�����(<�E1�����qr$�QVSI͝��5F�\��;RwK�2jG-��E��ڎ���*���(}vf%~���hHS�b};��ˉ ZJ=��J���x`��� /dȉ����v�ޖ~Z�VK����?:�Ϙn_z#0�����=jk�9���z3�u�O�8�cQO1�b�C��;F�����B���20��>3���g���X>"�!X�}t"����S�X~|�����m����툄�����m��!����=1�O]q	�!=�u ��':�in(a�
 L�g�M�S|�O��}o �W�Q��e!O���8���?7��\#K�AMo����ۋz8��������o����ň@�罔�|2k[�ʅI��|w�b�-N���6�d7^�K��d4*�
�" m4���x۲!_���bx����Y�^�rx����%��� ��':נ��I+lq���w�q�������ԙ���֑��͜l[�}�V;��e'm���;���W�|N����h�f�Tu���0Z�˜Oe#h���`�m�(�[��[{�wCi_����]Ʉ+|����(T��<q���I��y�Ŭ�x�r�e�}{+\L٬�N�,q��T�қ �r��oT�^�Td,�sB/�S,,%���r���;\"��',5�h���X]g*��y
�	�o���0�tWB�x�jOɍ���Z0:�!t�߉PW�C3��nH�7貹&Q��ʽ�3��V4����xӜ�:�:��bRȨ��gc�@��O�[\�/ADo�?�@7Y�)3� ��R�#]��[2�c��D��S�k�~�#�7@�a�Ӎ����N&ب
���R䂐3 ��C��ъX���(E��ټ�p�+;�N�w	�i��]K�4R��ceM�����-~�8�b���M�=�miS���IB"9�<�c�X�s�zS��a@�>�_3�W���R��\9�s�9D`8U7���/N��M5yՊtհdM�g���2�$����+�<�vO��T�ἠ��;:<���UrV]�~���~�r]b�.�r�(S�Q"NJS����!xjC*�!1Y1���D�q��C��;������e�������#mS�ј�\MJ� ���Mi�|�c��`�J���u�$9Kt�'��j��iI��<ǵ�34��4�'hG��?:�w����l�N4�;��dw	�Cr"xd[�{��!�]�?��X�ˤ��Y��gF�sO޾�K�ڬy9�av��t[
0ist���Z��GQ �p�߭��+qN��u����f��)j'
V[nD��Zh'�SASV\b@�B���k�J���빕�eK�z��f���\sᎭ=�=O������r�%j�^/r���6��N��E`�?В�ɫ0�7�9N��9FgL�J�"}�X�12�
/W��BzjzMT�D�z��x_�^���(Ū]��xJm\���s螺@{��o�^��!��Fr)��j7%�y����x���k��I�_����ʥ4�G�;�DK8@����hOb�l�3.�n����_d<�i�R-�`�R?J�����uﷸ[���-H���iIq3�.a�"�4)�9�������vx�y�	dg��G�A>��<�GRO���D���Uc�-�T�Q��,�P>�q�,r�T���l}5�9��c`e�V��"z����AC-�5��C���0��{�ʶǷ�>��?�d�B ��G[���y9`�����}׺���m$NۢW�������������!-�l�%���ݬ��[�҃�-�m���7q�VR��gl\Wv�{xp�i����y#��xm gO��5�Δ���_���>;[���vI���/婫����@�0��Db��#<3I��p�Qy��B�)���M�^\u$����t&i�瘴�ӕ�I���z8s>9�{4(�"�[���KA���8���C����6$�j�#��C��@v�^���AV��X�=c@71Q��26A�hD�T����=�_��l��O��������j�{
��������;% ����&\I-��8�J�ٲ��Jb�k �_�����l�������]m�ݾ�<+ݭ��e����K9wq�ܥs��w�Q��:��-�ӿ6Dt{�(�4{�L�c���Ř����H�,]�ޢ��2����a��y(��oS_:yr
��1�K��rL��1��n��*|*�
�
h?�7.�CV'�{�iW�j�@bj���8D����������{��W_8����.ͪ-�ԏ�vu�j�{�̫�'P�΄UȢ�U'���/F�m�]�`MwY�*��p�y�{|��oS��f�%�4�93�|.]���i����U�rXe�-O�2����^O#ʦ�=����K��]��D�Z�B
�D�KV�9�r~�5_	��^�=w�u�5�pʅ`|:
�cÙ����i�%�z|�(L�AW �=��8��p8�6o�;K6������ʰ��H��!V��l�×I[���P?cٷ���QJ]H�
��Se�lru% ,MWʪ�*�{�9vd�]�f���a�w� 푩��s]#Pf�����������n��k�bQp���ė��N���&s�q�hl��޴��lN��%��Frm��'�S�I��8Pmֱ7^��
�}�?�<�;���n�n�G�����<8	���d�[�E�H��x�ۨMSˤ5ݷ�D>t#�ʫ�B�pʨa���.��F�O�VՆ�f?��l�1���b2�O��q��	d���(��zRp/N�0�a.!`��l��RW��h�wY�֎o��V����_{Bt0��H��t���hC���v�6l<$WWP:UB�$o����qyVb�TO�8�W�$&8����IE���t��S2J�ɮ~U� �&��$���w�a�Jyߑ2#�<�|y̙й�ܼ���^"]�]�a��kr�p:�@͙~��ʥk�X@�C77(�C66�5��a�?�W��iԤ��"C෨�@��=2C�0�,��Ij���u����8ܞ%V�5��Y� #[N�Yf�P8$]�$tp�g�ӥx�_S�-v+Ý�.�i
nk�KK����l�Vw�0^R)Q�~l��d�9� �b˨k�W���٫�ŋp��cW�����c���v�����̗ɲ��w�<R�Kr�ɜYin�*5��SM���98������Ƽ���x���8�@</���5�\��b�8N�o��qC����k�v����R�Y�����TF�"�ҡg��ON�vO�D��y[��d�tч�[�*5]:�v����|�,Ig �jԄ!^��)�z{;E�9��C*���KKW��F	�Ol��&�;[��v�#�=`���oc���6Mijcn�y����ٿ��Mb6&j��"�I�@�=d���qh'j�4]CR�ן6����Qʃ�f�6�e��:�R�+Ξ!��~��)�%yJ�̄��2I�0�JS�f�f1(� a ��5�I������%3:ơKV�X����TAB߫��"�)��;�^��G$XRE��Д.�����$�R[ϗ�#�!�aq��4W��Ȑ�P}�Ņ.iK7n��,;�����TE��/��ϼ�#6�gz/ࢃ��
���Z�]���î~)'2�}%�($���+�1�����#����x0�ܵ��h���*Wi��`-O�=�jcz+��;��Z��x�WHI>�ȭ%*x�D	.���	'��Z�m��\�\�&�To�6�ѻ���Da�>rq�2�e�~�3��bH/2[����zu��s*W�/��|;���H�?�h]U�.v���$�*Uz1|Ś �9r�#'Q�'���6c�3��"�[���20�]T���e��[@����p.#�\��Tf4�0�Ԩ���7�B���H�w�n(r����h�Y�J7^��1\��R i��4aP�n���Yq�)Hp�u3���j�����Z�@ԕ  &�����x�`��w���󠂑P7�M��;-���S�Q/��>����enG�9�6���,&A��CCp�sG�緸����$W��r�}]}]o�#�z�39
P��3 j��h)E4�$8���^�7zPX�h�>�1�?��'�anᄋ$]��O+�(gp>5���-�,s���xi�hٯ�P�� ��v�}�Wdgk�s�K-�̜��.n��ll��rt��wl�`���1�����y��d滷Y��#�U?���ɧ�yG�i�l`��5��=jZ_�K�!�x�V8�>Xۖ�A
�q"�U�Ǒ��>�Y1 d{��:��#��mHq~&iN�~��8nJ�)��TlW��z�F�`��ʴq��?�#�^��\�KOy-7����PZʾ��^g�G��
:nZw�J���|�~3�t �ƀG}��Kq��ѣgq�X����;�A^�"q��-����=̔��1O�����8�,���ӉT`@ػ�/ζ���	R���P:0|���N$O�V�v�Af>�˚'m���ᝅ|¶��3�vF�-.�ޮ5u��E8���
��z��y�u����>�.?�4A$�N����y���cSy`��{Q��WYK����%"�m�� �cU@���,�rX���ϋ#}-D��1�>7?�EU��jG0��=���q�A�G��X�2�t?�`�{��Y�g�ƤS�\m� 	PO���u��A4���o���OїJ#7�D�u�~nO?�Σ��ާ�BQ�5rr�~��E���O����y�"�]F��e�_��_F�D�6k���>�ē� FsXg�H[Ǿ���ܶ���vΥ-�����	zk��C�P����M�PuB���9�/�C�@	@�0�/�M�����lu�d萝�h�3hҒ!͂[��9�@��*.d �u68����Q����������Y[����j����� ��@WE,���e�u�qvǔ��1fjM�N�Cq�ZQ��r��D�E�!��v�M��
����*�O]�� W$pG��4��#��څ+�Q�s�.��CD��b?���pg�#��� 	@���wU]@�t�>O]�yiĪJc��g]0)��a����:H�_�&e�K�����-'0\B�1�r�,t�6dcڅ�/�$$ )*g"�r_���W,!�����ҷ�FǺ9>n�]�l墍��Ƨ�`A��W�\���0篬:��:�T�:p��`#0�����c���;���b;��uL���q�Z���	�jp������Q�C��nq����ZH��I�y\�
�-�d�lW吡�?Q.����&Q1#�@���(�W(��B��Lײ�EW�x%)��_K���[�V�h�\BJĳU �Z���kdۗ:��ɡ�&���Y�gqcO*�<>q]�o$�]�8�]�������*�(Y�i.��yT�oV�Sa�6��;J�	�l�Q�g��%u�n鏙�N�Y�-�T��О�8ï�qyY�K�r:��n���F9Q��� �D$-�:��sEA���l��2�p\��h����Ys	�A�����|w�w���V+l�W�k���E�x�p�"C	;��[#j�.Ѧw�nQݾۡE*b>�m���M�㣍�]�P����"��[x|)>�vv�Ky�m2�����ɇ�B�#=���4�W�;:�κ��`Ւݽ�z�N�MuM�Q��,��0����V����)ȋ�R�`��O杆n��|9���$ ������آ�`(���@��R �1��$ÿ����j-��2i�쪼�v���D�L:s�[���S��V�����I�)ݸ�^N�dmfu2�L`�I�)l�����oز��p��a�n�۳K��Vo�������ۏNI�n����}{�tVc0�)�;�&�:]xA�qa��m�m����D�_
ūٟ-��1����w"�gk��V[u#?�j�3��F8�N�1( �>r�s���JS/d8i�I����ٖ�P���n��&O���q���ҧi(%����Cm۩�7D=��-��w�	R"e�Da�pKRbmm���]*wEt] ���Jk�Ȫ�}����KO����*���.�C8��C塒��k!��L�b[� �c����)c�b��xnz��h��_pϛ�v��'`)�Nu�Dw&�9���h�W��3��p�͍�(4�A��!v��|(m��z������6>.���c�e	\� Hc �N�>}�wG����d��"���DJ��gA�;�&i��B7=g�T��γb� �h�fN�_+��i4H�?R^ݮ.|�G4���9x-��4���	m�d�!0D��e��7U-̠J-����Xa�o��D�dTi�g���o�oeJ�yj�.'+�A�q���p�c`=�������Pw.@�SI��Cz0��F����DL��I^��=T9'���C��ė�B4�A�ٜ��k�fh�R�ÈWR�n ��8 �w�o��!Q�	r�*�jX�K���c�+K�������$��O��5�q�
�q\'��ĘA��t��y�>�ނN�3��NH`�9`���ӿ����M�����7������ۗm��$��ř�rWɋ�5��b"S��\�E׫ʸGB:T�_.5qC٭��R�%䔽��S��.�-I}&��CT�ڂ7���:�U�S�f�K��^���+�������ڔ~�A��g�N�L���=|}�� Zܰ��gx����K  A䈿+�A%yE��(�kӞ���fI�a�tHzO�^�<eڢ�M���@F���@���$�Z9�����w�@^[K��R�k������e�fΞ��7�$=���˘�-s�b��p������X�l3m1z��P$��ʔ}6Q�-����{_�'����Sx,bG��#��g:a�W[3�&�FӐ1&W�]�T�	@$v{0� zd���Q��77h���g9��&�����>��Ũ��C���0��i�U��r�N�M�$Ċ�E^��5y�a|�d�[a	|��Ȃ�qDx������N�9ōIރ�V�-���[*"�O��b�H���@9
��v7�ݼ)X0�\6��,�V�Z���w�6������eĬcM��+ ЗL]$}�z]��(\���xk��|rb*���}Ć��؃v͇R	-;fc�ߟ[U~L �A^����:H�i�ϖ�2��b�/T���;	����G�sEv��2�=��� �Y�O�1�����Uw�S�U��Y� �i�6n1�)W���������e<!��U@&�.�I��5P'�5���.N�+�[�+'�g���R��V4e�:1\^�sp^s�e�޲X9w��\�������
a���U��nV��g7Ѡ�J�*|Ik�����,���Y�Ǵ�ғ�V����BQ�Z���z"�*�l�3���'D&�Y�eei��&e�5�8F�o���[��a)�RR��ՠm\q�b&{@h=�髼�/WB�ѫ�}NH��ټ�T� �}M�nz!$|/��M�gה��?Q&���Y��m`���N�Yh�����g��e12�<q"�P��7U�T�ʄ9v��=@#�Ӛ�����a
��c�-�Au7����l#|�Ww��?' �}� .��� /�~Ƅ`��3��+S�[q�:i���3�f���0F��#}�Ѡ�퇦��&��sh�L*�tKЀ�9`��]f�!I�s�V�oX^Y���~0I��?'��ZUp7���I�}�A��ئ�Q��
;���ܪ��	4�����Q�c�N6I+�!��͍u��g>^�� ���'� �6���w��~��<�z���ghk6'�e�+H�΅h&�Uҽ+����.��Z��.{�:Aj��f�!�ډ�j���f�^Ȁ�"�x6�Ѳ6�^:�|�n���PBo>�9��tM2�
��uM12�A�#uL�M�\yCg��>p�~a��ˣ���pt �m����=L�9~�p�*t��Eq4H�Ut��O��X���~�EgJ�Z��s�3/���wHZ���_b�#��_�[�%�H�O*@��4d�8���Ș�v@=��j�	A������zT���l�~
�p8��N�������!!\�rPP��Ӣ��k,t�������2�*��8Ԭ���؇iR+g
c����%����&�P� a!��s�YtX�^iJy$8���g94DU��B� �����p���՞�ʈ�P��E��k������.zdf tw״�?Yo�pZAgzbj��P�����wsJ;@�byLCn�) ���[���d�J'��և���CJ�������"LkזUuL ��߰C�tR�m-���T=ƗUTsJ>�ėA�������Qxj�MOtaH�?g���]�Jd��	w��]�� x�����L�(�|pv@��bu~	Uj�o��:2�@(�*T����f��^�&+cQ�S<�� ����M�Dq�&h4����vT+z0dڬ��� �zu7cv����.����^M�Q [(� ���4��},�i9�+��_�}�I����Y��!E=x檶���2���@�?o�BR�/�^�VR��#�xk�M.=�t:��9�s�u�O�	;�8Dv}fO5��wQő��jT�)�-���G�A�?�2z�"p�B��9f�G�t�� 6	���ӎ�c.z��I~���#�+�{~�1�i�9Ay���i	So+=�z��W��i�(f4�-\u0�	V���D��˿Wl�՘F�����N�=p��Z�⬞�J/��(������P`�� �+ga,�c�G�����T����ݵ�74�|ϰ��6��ޛ��xH�]ȇ�G%&����;#F�A
t����y���?�Ul�����\��D�E.d�e�p������g���y�n3e^_�ɵ?�2��s�jɿ��ub,\��S���r]5�X�|6 ��c�C��U\�m�� �:���'^l���Ζt����R�nZ0P/_����XT�m�iD:���v����=��R"�6������-��)��*��B���yS��1&�I��w�Ż��yS��A>�yU�w�&��1}�w����D�G���ԍqfȌ�6��m���؊�iC��� *PQ�$����@��(/s��qIb�6U}}g&�P��u.��HP���(a�ZԒA��Ô�L�:�lF��цL�K��F���hv���-�^�F���#f����� �1Ħ�v�����T�2	����x��W�]��Qh?��!�v�ӎ��^U16D︧}���Ve\�q��Os�~G�q�&Yɂ�1 �� A
:��p<��"կ>�yR�=�4"�����<%
��ځMO��t�D�h��~$2�ceɟ%����(@��/���@��֟D���hx;�D����Φ�����qz�g+���1}8�lc���z���V��b&��,5;�{�Z.��6� ��	��#�S!5t�=2S�t7c���b������0����ɽ��z�G%�k��w�;���u�	���y�ED��N|��\���f\���� ��l�gK�t4��݆}���4�OK���
Xe�V�Ȯ�7Jӓ����L�q��WJ��7�8|��!:�`)�Y�-��Pa��
�X�8eτ������5�^�Qc�!4H'�=J�?������0{�=>�l2?�Q�+�tbX5�{[�cϢ�]u�'�7��K��*b�v��f\J�mdkũ��C�O���R���Ei�ێ��C$Ng�՘d+��]�juÕP)�o�(�S�
���N�{�la�]�Uشx�.�������'l�3�q� �W�D�X��챪��Kz�8m���܈v�ĳA��MP�V�d��Z:C��#ݿ����Z�m5S,{Q���C!����cX*�D�!�^�i~�W�-ZB�bH嵌��xm�:��S�a�f'��L�Kq�_�DrN2�o��*��<7�F��av���o����-�X���y��az�JZA���j���5����9<E�����O��q�¬��c�L@�|��ה�h%�R��n����2��6��;��퐺P�96�&�<��W��O�SX����������0߬ 7!�X+Nf�:��a	����#�g ]k�Ҩc�j������OG�p��_�Jo���n�k'�1M��d�7��S �%_�*80����Ud�;�6�WAi(w��M�5 #�����*�H�"jo�����Eyc�U?�)��b�y��e�=mNaJ̵\��Vb6ɿR1�M�$TwyU�����'C��k��yE_��/{�q�f�����1��P&$�ŧF�l�H�Yo��}�7xS6�]�x�h�n��A@�Y��y�[,��;��Zߠl�Iˊ9�eWG�j(���,QT2Q*��M�_����~T]09�|۩��R�A��M@��� �x?�C��Em���*���t� ��œ�V=�a4�'>�*oN�(�}ΗJ�kY*��$��ܓ0+$�9N�����z�C����:�cS.V>��F�jg�ﶣHF|�@�=�Kb�v[蹞 b��`/T�)`�X��|�Ȉh���O[�2�{��:�p��m��qL	�eix%A'lS� 	6v�n�"9�-a�M>�VH\�k����N��!]]�uD�/|��/(��zV��*BQ��p"�fG��Ε�;.<�^�	���#ap�Hrg��d��,
'���\I�k��
�f�_�Ĺo���c�R8`�0�i�Z3͑�ЧV�H��2��P4O�mr���E~���h��:��"c�~��(�����I5�5>��$�>>
��V�փ�����κ�ű7�������:)��g�2�{�̳���QS���}A�98�h:�\��D@U�T�ƴNS�8F����Z\�7�Bd��Y#�f�7�p3(����	�X��@
Bz3c��Nˣ�b?_ЇmC�Y�F��$8���q�+��F?7�"�e�@P�����yvv��e�5�߫D�+#���3&츁���0)�8H�Ҳ�R�q�7AN�K��Į�Ny���2�(G�0Kod�&�G�'#k|�ð���%���D�� ��%7��/�+1�B�I��u��d��S����YV�3�����O ���sT*���Ԉ6�ΦW��7��k�%�#*}�|/�:蔦0��Z�!�]R/��� ���;����.?6%�,{cf$�y�V�@Wy������Z� �Ǥ:�Ѐ�q�ᙳ�**+@�90ד �V��R�фf��,�=� 1�in7��rg�:���c*��Zm'�v��uw�T����P� 1�D��)�E�+�Pp���	/��H����]��H���|�0V܍��<��t�m7p���0Xt2��Wt⩀@�9c�ζ,��;*eGۑ�4c�ʙ����o�=�9�<�������q�d��e��[8�L�w���z!�2��c	��v�\.٣`h��-����!ũ��%�r/YL��_�L)�~V������%�ȹ�����p��O�kh@�n��m[�koW�,O��Ό&1g���.K5|�pn�.�wk_T���KG�Ѝ� �*��=O��g�[=�
LE�nb���쑼s���ǝ�.;�͹6�0���1:��Z~²�ҵPld��Ӵ_�Q�^7��7B�Q�KT�E$&\Tb�;*s�fw�ݵo����4�(6vG���b5y{5@�|���,B��ڴ��x���K��w��.��	�pn����V�s��}I8��:�sI��&�?���0U�h)	�����K�ᐚ����cB���&cO%
OCM����X

��A�,U��]I<�����[���1����@�-�`�*'(h�u��"�x ��(�"s��� �4�۽��[U<*�Ϛ$w�Ų-��v�����Dˡ�I=&x�R��y����c	Xp�����5y�	��T���ۼU8���D奾z�7�~/,9��*)�k���_߶��B��R�0j��e+��q��B���pHKNBKxN� ��G�y\2<�P�x"O���N����ym����'F �� ��B���g������!�Cw&���X[Yɸ�����e�=��e�1p��hE�bf�j��M�
�����G-?3��� c�C���5R����D6?�� q�`�&7,|�ZB��-� #�s���P��%#C�c>ew{X(�F�8���j���&�6�m'9��P��r�~Ė�CoYbS<q@��]����c��с2+}�G����ޫ؝��S�T���x�����Q)ln&U�F�t���LwND��Έ�ჲ1 �29���A���9�f[
B;/Y�r�#U�vpE�[���Ltc�uy�h�WiO��^@U��������)C�0i�&)D�K#�������h�8��������h���2�_��_ݱ�ej��;�{�+W@C���qx���8���F�/j��sgUw�3� ���� �y+��2�WM���U���4D��YГm�*@�<3sUB���{Pׇ
Nh=,{�ՒM�Y���m%��c��ˮ�P��t��h�z,���z�Ő;���[q&��M�A�8(��e	��J�A7�)����E�j�I��0j���M�/�Ɍ��,@X��I�T���ćU��Zj�k��H��u�+��4"�H$y
+�^��|��{q�ܰd�c�Sz����A�Cl�M m����?9��=�u�����5G��W�%8Y\B�}B��r�d[�����j^�+p���u�L1tw��-�M��`g��~R�݈�^���R�c�X��|�
a5Ǉ\4�F�A�5j�������4�X�_�J���Fa0�n�R �J�w�Ѵ}�IN�Aط̣w!����pcO��ŧ�rҁ`<�ݗ���A��������ҟ۽�5
o��4DA��ΰd��X���XU~��na�C$'-&�6<z�K%1�a�Ҁ{s"RH_'ĸ��)j/<��v9�#~��nT6��Nd;N+БRfM΅|uy�E��jC׃�����_�,Q���:_���S`�p9`n�?��PL y�Jk2y}�40vV�H���>t;�Hf��w���[�o>"��Դ�*�1�+��u�M��,��~�H؈�:�ޛ�����AA���˛ �lp䭷C��>w���I��@�#j٠��'{Kц�a����I�s��"͕K�iJ$�p�l�/Nd�1D)��/i��=aO^�T����B5�Z#B�ǯ�Y�S��޳(�	�d�}����#,Z��bO�}��a��R&�����04�.cʺA��Q�L�YX_��[��߁R}�ɧpA^�`�������v3���{W�N<��]��9���8H��"��z��r-�XLZ,����؋��M"�E�j�����5��V��� �2I����T`'7�,b�vC�����d+K��b����B݋?{���q�N�؎M����dUPv�󢀔2(��͐���ch��o����<n�|�����􃎕 M�����ٲ���d��tH�z\��@1�P�~#��Gb��t���T�"cے�5��l7p���g�/ڒ�`�FP	�I���tS#t�6����K%��.�F��$;��żD��
52u�u4��(V����(�+=�J����ws3�3�����v�����c۝�ͻy4�"�<zF7�0�H����fE� 0
|���7�S=�]'�R����CH�?��Ɉ9-!����v�FH����h�P;��M�}TO;�3/�dw_+Ջr���q�VC����0SD
Cv�ؽ9�B��Mʬ��S�Y߂	�� ��r�j6b�-�xL�� i;��0W�)��h�~�2[�!\Βa��2]��D�� ����z���H����>���j��uE���|�#X_���`��k��$�����Z]ӥ�Ԅ���tt%wzEX,���	I�<�J+��]]y��"���L+��i��R	!���
��ؕ�A����ɢ�>*�����,g���r�&Oۧ�e���~X�Ie��g�'S�(��y-�y&2t舤w�B�w�23��c����P�81��e�A��=�?�&p	1ZC������>R��p����@E�^/X�� ���'k�X�B� �?�$y��j:�}��}���<�Z�Ʈ��1�������ʧi;�?����%k���27��=��ta��b�h�\b�k�p�;��GU�3��Y���`b��E�8DPNݹτ�S�[q[
�-k S�Je�q01�_��M�L�v�:;Q��/�u1K�A.O�(a�sd�+c����ٓ�=J��ѹI�b��l�_���]����W�5|MP�{Ҍ��v QՍ�]�Mϊ���r�����2�Uw<O�ڨ�+s��uAm�{����<X�T!Z�V3#�BC��S"��i���w\�W�0j�;j�F}�o���F�8��K $v��1����92�n�'.�D!Q���+��ڎk� �fK�
$��d�Cɘkꛢ��S��U����N�X����� �>�j^9QɻF�B@�wG�(n�J���׉�TfŕO��n���d��^e���?�F�xLT�Gh
*�B��qԨ¦��x?���`;/~�fE/A@ď��o;�1E�� �!�
x���`W�66�_�����GI <*)�$�Ij��s��U{,��Jp�{Ɣ��#%��j�ް{d�T�H�2�N8��Ё��@�v��0��3������P�#�g�z;���zO�l��f�(��+f�s)��.������HZ`����N����
�˞d���	@���Y�8��L���(hSD@�UH�-�w��F�U�*�#n{O�a��N�kR~�D礬ZkQK�V&��/@ͻ����p7��:��5�������7[=M����*����5��e�\��ǤаA9�;�	�
��l�n�Pao�ٕ��72'�s�����Cz��������c�%��!�H�/6?K��%��L�r^L�b��f�:�X��y|
�i����h�N�*_5���	5-�X�a��ʭÇ��,!݊��d�8��(@���1�c:����v��)�P�-�	��S��kPs5�9!�M ��Z���9��w��ttP�����C�n�O�{�*x�sU̇J����xÁU�����ɄY:��C����Ix�Ԁ��
�׷\B)%�ф����k�x�g;���uP�k�m���P�mz�x_���$M|jU)�+�&����J	MS�Sʓq,�g��& �ϳ���r]��IJ*4�G�ZTG�֙�����q���\#���vE[��ݑ�4���Ȯ�^�� �:7$]��y������O�|䍧���&��Lk�<tB�D���!�,��q�"�ʈ�T9{hr`,ՙ���G���w��3-_�^��6�B�a�Ĝ�d���V�v]����m��rC��/�n>-���k���1��~�_VH;�6�i^ƽӇ����ΰ��P��Z��~O�-����Iu�y�����/��S��J�2Q�k�*@�b���7R��в��]ܒ0`x�uyq�3���G����|�E-y�F��Ifh��ۢ��\��F��r��p�!�
~� ���x�3Иzd ?y�9�A�ɀ�=IAXgM�ܨ3=��嘈��Q�HX�`l��U#����4d25�����|��ٌ�nż�]���&�9=Y�B�C�/H��-�ڀR����m�I@�ם !��V,ʑ�"%���Hz��Eި�$�̢ Q�/���D6i�d�Yݽ�f�g�'q�w�������k��nO\7�T2�/yX.i��j�����J}��������j�PkT�T\��.�S(l�[�U!����	�Ony���Š,��pH�#�;��[�&�i�'5��2��t��%����g����M�����{j����'��\����+ ��i���Ě]�*�,t2���<����"�f�TPa��~j[�~��Z�����3]�c ]K�~
H��R"+���}l�Ze�л�{	�:���M3�~a�Bf�p�)KP�] �3u�f�Ӑ5��X�<���`�k��#����}����Aqc��b�����,��S��ؙ���
Yqgc��$�Fj$�"�S�wƨ�םe�R�#�8w�sk�5�v�mz�b�,��5�}���p���&1S�o���E�~�E��E�oyP��y�%կ$<-��}�Ҫ������$��3��95�sQ[�!>Y~��+r���Ty�]�"~�b����<��̡Ԅl��DL)���J�7*nڡ$���YMX�W�02��rG����e垍'OPZ��������ʮ�1�>ܔ$K�����Fj��̮x4?�����J�-ZR��7vܚl�Q�SH:]9C��iGG��0;�b�y���J�9��,zL�ˍ�����u� �7R��#��H.�7��̩�Ձ	}L��z����?]� �W��hS������f���|�9�M��N�!�	��2z:exl������lxng��2����^�b=հ�.ꩿjr�>WW�|6��e9|U�>��3Ȟ8�2+��Ք}y�p{̕2IRFpĲӳ����������dw�ÿ��-/ry& �z���؟!l�����hܨ&fP��1�"�T�$�S۳�G�vZ0��eI����X̵1�;�X�l�0Zo�qr{y}�Y˔��(Gk��0���׎�;�%Uˆ[`@R�n"�[��qH���"v���~":�ku�11�����p�KT� �q�X c���2��>Oܹ��hĽ�]߆��ƈbQ����.\�ȊHQ�==�y�cEC<��{ʰ���o�����c�6J2��������Ր��N���!��+�c�:KeޝgY��q�wp�`�GHeD"r��8\��&������,9s�U�J��pM�:�����mjys	���������e �4Z��%�G���\ G 
ӽ�gR>�Z=�ۉ�����W��`j&!�C���\�=�|y3�#ܻ~��;GVlU;q�2��K����,��t*�5Ud���b�*�6͹���r�ԈiG�/�zT�-���M�:�yk�<��#St$S�!>��q�� w��U��
�u�w~�֍�A�:z�#l��
�~��ڧ^*��)���\�.���� G⊲�p�Q��Y=�@��{�����`��6���F��1�W��n���+߀Ո����]�����%)�c��Ofd~�X����~T� T�n!�{�,��d,]��Ux�W�'a^F��R�������{��R��=?��H�a��T���)�g���qz��"�Z������;�+�^�@��dJg��!e�+)��(r�f(E��ba�O��$�F��u�cڦ)�ȃ��H*Q-OuźH�z�����!���"����n��8-� �|�s�ݚ�p��0�_���W�oq���`k�M���X��E�z�#&_�r�2t��@�8l�0d����Ψ0�oV�2�@c�RF-�p�YQ�p@{/�7Ej���&ʅ���6r��������b����� �49��X��ldO�{��R@	|Q�"��S5t��
o 9�L�z{B�������U�$�1Ӝ�$��Lk���\���5�Иl�?�b.�6��S�kk5Q��T�j |Kh���) ��NvT��XV�џ�,0��Ox�p.z���p�S\v ���L#�6YE4O�ӛ���s�m�ۂ���9���}�u�����~n�y�6$Y�t�iN���$۩�D�_������K��\5���ʬd	�!%��������P���`4��,���.ߙᑨ�&�� M(��rt;��V�VR�.t���ΓŸs;��Z�����
%{R�dIj��E�[@nJ�>޷5縷�J/��<l�f�h���~���Er��b,�(tL�P\&,���o� ��{�c�iJ-l��K����!:���<l�����Yz_Vi2�$B[��y����{<�Y���������ݺ"#]�`�׳S�3�|C�3���C:93u!� 3����rp���5ؾ hp˙fXzi6��C��ץ�� J�#�r�D!��ؑ@ ��=���/��cL���/�k�4,
�5�1� E�U5��$O�^`[�𓆵S�X�v8����G.���E ����ȉ���zLנ�"O�)aP�r#�;W��$�s"+]LkZ0�� �L�$����S���9��҅�n-؄���M`�&�N	�[�rS��[۠�y���P̼+�~:*��X��@\����))9�  ��|��������Ɛ�#R���M((\�3唢�
bcL�fz�(��Q��rJmU�qu4�rb�#�PM��b'`�����F�+G�e�����D��)«:��#p��Y�ݭ������n`;4�����Q���tƉ+B����K�G��Q���F+#�9��W�7���,�Sg��o�O� m훮^�O�l�紪a�o�Y�q����#d@}G��:(��z�`>N`�/,�+��;5	<����i�a8YI�G ��{N Ui��ل�Y�c�j�d=��Ԡ��z]͑+.O�r��PiHӧ���Lr�^1�aTjoX�%�	Ln�ˡ�ɯR���A��9�,Е�ee��ΖL��I�W�h[�Ar��L�,�C	ҮK?'§�%����|�d��a�_���º(�2鵧c�bq9�&9q�[�7�w;:4;2�c���?��Hr��A�*I7�qU.�-���x�K�E���������2~�F��n8�e2�ۃ�̆�Uh*��
/��@�tX��قى��ҧF98XI��!f����3sk�#�cCc�D=_�Hr��a�K���t�p�[)�1��ΰ��yvS�D�x9�bz>��l���ѵ�ͼ�[����0����3^"^�9m�����Y?q�]…�A�eC���4���t�0̒tBW\,�sY��ϮƉ;$�"��6,�X%���9�g�*��W������%�D�혔��pd
��C�%�߶�5��`ъ�<h恰�yn�6M��h\����^��*u[�M7�:�l�.�ϠQ�u//>s������
'��j�R��%ɽ�t�[��+Gry�$U�0!�80�,ē<(񾧀Fҳ��|�찍�a%wh�3R�0�v���k1�Ι+8�M%ԛ�|��O�%�t�2�EB�oޢ?���p:��9�1��_t�?o�d+q8�ũ ܓ��!���$B�>�1:9g�?�w��zk>�?��$pH�<2�3 ��|'8��=�\��D��1̆XW�G��ί�˙p����`��֑b�=Щ�G��b_zj���w&�ч����������:EW5��Ljq�\�[�F����f�R�b�xRp��|�������j|��g��K�v$�,_��=�)ы�Wþ6�?���鰃�K��A�HW�遮4Lɷ�ح}����je� �)���S)!)����E�}ms�̹����0�{�3���I�
lϴdm,�f���2;I�v~TF@��`'��	���AơBNhA�BӋl�v�/�T�+�V�h�k~fV��aē�IZ$�浙H�1\��]BC�[ſH�k�9�`����a�����9K� fGi��du���aL���vo�;P����ĐI#�%��4� ����_�:��+��R��K��k0����pC�2F�GRW�u�_��$����`@�߭��a�6պ�cJt�
;��(��`�B}�'�m�=�aP�]!�tP�B��%!��}xr\��'F��]@���u<���=�#A�+=��_�B6H���P��
v����ޅ����u�H�j�i�O���|�����UoԶiu�`��V���|�.�%�^N	��6�<�T!�̍��M��'�TÁ7�H���#`�����X0�!O�'];�[�pW���{lV�"6�8X:v7�be��x�+zTK�n*y�9އHL�(;���2 _��5F�����������X^��o�]�P.�A<��i3��PMzYWI���˿��y�ə\f���U\+a�9,"׌K���7���[e�،�ny2��M0�Zr�R�]�}:�&�kaA}}�}p��ў�O��4B�d,Z؝�O�R-9$y�L�2D���P���G*��rVY��>�[b��l��a�i�b�r1�S�eqݚ�E�����S� +(e�PZ�l-�n��][���,� �F11)�bD��\Dv���q����x������î���c+�M(�tS�l�K�-^�@��JC�����O6���r𦆘){�'�e����7_���_���i�0��5����-�h���fܻ��TYh�,_Ҕ�m��q�S�m���
��t�U
䆲��������'h���3�/F�}�quی'�J�^*�D�;�ÄYQ�0�Z߉��)0$�Y%v���WF��ٳ�ݓ�n�� J���k�J=i[�jn�'|W�AE3�g<+��R��V����fJ��T�$�g�������a���ɠ�Zro�o��b�1_C�I��C�q�p���^*N6�\Mvԉ����s��A��+o@݌����﹨��#�D|f�Q����R� &��g���bQ?���J@��f"���}��ξr���U�:#��k�*T�+YY/ GGRJ��
u;Ψ�z͸/
����7�1ߣ��:�-��N^�cy2�֚m��!.\�ԟlו��Cʛ�رJ���io���@���*� a��H�^k�Ԡ{�~y"��ts�U����<S�i�g��Hx���˼y�O��1"�3%�x�ﲝ��y:4J��\��h �m�|�@@J�+5�Y�h��a�gV���ޙ �D \���<��I��$_��V�w����������n���V����s��#NE��W��ͯm�k�S82eBr�b@5���6B��y��%Ŕ,T���BDO:�X� ��7��ۦ7�6��H��� � $��u��7�����F�EUW�'�5�n��)�{m���4`���
�7V�,��ȾM�zEhD4�+���F[3�� ���q���"	�0��`j���� ������ ����H��
e�Z��1�%���7�&���˕�Y��������CW�L�0���	vd�6:�V�3'�52��Z�d�7����it��(Bq�Gv�����ș���|��Q3�[>c��@��@@z/N����g܂�����T��)B!��W�3�F��ea!�����ɫ<w�1U�.2��O2�\��A;\�<�T�r�rg��Vi*(�b�������f���b�6�|%H��!7w��)�X�0S����n~�p
���&9g�{ͽ)m76�L�>�x
�7�2wcݩ�n�]�)'�''�h}
�g��$�t���㓟��
��B���C��t�9ĸ��b���3����	"���[�)��h�M��J�����L�Q�:~��gU<8J�=�_F�1��QrIL҇A�-�����	u��տr�f�D	s+5Ʈķ2�������Nqi�p�摀��\��n��L�U tt[+ў��jM ����I���.S^ALǙ#G���z�<�Dxf���W��˿�s��@�%9�]IgЍ�֠��n덅�ɝF;bHG���Y��-��S�vR�,��Յ�fE��J�1mRH�{��A��̷����mrkh�&�Ii�ovXd�O�JU;��e�\
1p����� 7�j���'x�0�r��,�}ߔ+��L`TG�J�X�3���8(P��>v=�i��z#���$����Hɵ��cg��;�0S��ջ�����t�i�7|�	v�`y+��_ %�{�"҉%8��H���kA����x�� �G
3]�]�Q�S񋡧��S���)��������#�.���CX~�����⡬X,��)T��3�f�P�.����V��.
��ҊY��^>�e���:����"ci�9G4�:�+q�-�ަ�C3��AM�r���)F� )^�:���i�Z�u�^@?&^���d�/
j���D�1�baS1@$�Iz�Pe�|�&Q�g�� �Mo8��lj��Ḇ{۴<P���J/a��>Am�b�Fm��6q�H+y���=Q��N�V���.�L*���p�)�E�Ɵ�2�G-9U��̅P���J��
�d�Ux8����r���!4���q��h��e�������U�F���m�7
��d�<+k�>�nt*j8�g,��Erz�Z�1���y�h0><�`�	S�.�����+>�+,��;��MK��*]��Ÿ�	�h�'~QˤK��a����{٦�.��XS4w\���#l�@�\(:���v�vH���0�O��K;a#��N�O��T�B��^c����x����GN喞�,���h��|�����o-�'|���ϼx��1Zoa�_�N��;!��:�=�^�',�`�j�0=9Z^��}(�_?�r�����CYT�D���$�!ً�,���
�~)Mi�{X%����y��K�a�8����K�]Ć#1��B${Z}���lx�=�u�6Z�k�{�� ۟��i����Y�)�P��4+�*$��o<��r�����<c~�hL�y&�ʝt��B-���K�ǰ(��H�/b�G(I�>�m̀�y�<��X�͂�3c]�Q%5����U=e��E\���C��������Kѱ����Mk�^$���9]��Q|JAN� ��G���&�Rw#���JtƯ�rQ��'��2ˣ.??��<�xf��B�GZaӧѢF>��*��SQ�	�#�mr\�H��Ny+�f��4i܆�tb��I��G-�
��-�]B��.�2�}.꧖��j��Yd�F�N�bHD��`|�f��E5#8K\r {����]���Im�o_�g9w�B2}{?��|f���H�v�O<��Um�k����W��G�a�C����x����oø|�V������X����ߨ���Q�}�ltv)�ϵ���̀�A�y��ҡy��VW���v���=����h&��6U���&ϒs����z�����H�2�?�&!����p�&G����I?�#i{�]��?͠��,�[*f4��=rAjY���-�b5Ґa�o�;��ш��ԡ!M�Mr�p�c�0ii5�=?2�W�=�2�#�Xؤ�H&�p�a�G�d,O�];F��}���p��P�_s��oV��W�Cjw�eА3n�%l�N�V��_���pdj�2������Df���kU��$ޠV���e��8N�r��_���@��&{���y���v"�-e0���Q��T�"Bt.ϙ�vX�#O%�����U�	c>��JD�\M�$PZu	Fm%�%�8�U�X��ڮ20d��|"�zo&h�"�q�<�=y�vFy��M��L��F|vW�`�����$�G�������h��-un�n��2@f�~�u��uc�g-���"م���2Z�t
߳�z��ff؛D �F�fw|b�K�rCV����V}+�\�_�����"�-|PW�\�Ȃ7wi��Ȥ��	N{#�)C�BW5�i���7*~�2�cj�#� ��Uf�5�g9��Yż�]�mud�>TQW��X�gƚ3�muw��i0�����m��
gR3x�����,��v�n%C6ei��A@'��!C��)���Μ},�?�p��a[VA��~s�R\��v[p`|�9�`�e�q=`�7�떡�_�CK��9�>��u���oSeWQH���%�/�^�����U�B�����e�c���ǘ'�`��|r!����5��K��"��:/e��T��)����@�"	Ԙ"sx�PM�I�`ۺ��ß�:9��T�!��8�ۉLtX��'2��V�N*�Z���c�6���:�B�Q	M߃�I�S��iH��[a: ��H�ʉ���LLHf�yqݧٷ����E�3���C�L��i$)����I̫��=ݔy���m�̿ia\tS����8E���q&�-������K^��ԣ��)�D�E� �wy�Lzꀩze]QO=H��|���l���	�bЇ�rg�-��������e����"�<�k��傍���r�P��D¯�3���h3{��U��Ϣ��k��?����{��B�e��Q,:Ω�n$�-\��G�����HFq\}�/$?�<�������۩�%#��8η|��Ѵ��}ѓw ~0q������&x��ޟ|��K���sj��4  d7�f�R�r�_����]M��=��P���H86,�{q 
`IY9�!��U7�,w&�lJ�E")���ǁ�����0{z�Y~4�v2��íݜb�Nm�jY��	X�9��0��e�?��{H�x7��E}�l$�V��N�qg����V�w�����V�����l7ów:j��!��C��O\7Q1#C�g�)���IA�P{�Y>ֹ3O�Z����VC�7��76!���,���߭��AM��sg��etj��o;��X���t��=��ϡ,�<)_�k�4?��m`�Ric>w��"���\�4������T��!�{�<f��z�[[�"Lr1�A4|�J�;M��vZ�_���������.i�� �|���pP� u�_�#�`.9R�~�Z�׽����O� {-�HG)��v~3���%h\�$���r%a� ��y�A��O�F�c�C��?�a''�i������J�9="�@���2�;��"�_#R~���+�tDW��S�s*3=(0?���+1N.�0��@��3d�����E��6��yFʱ*�,�S�p���1ɣ_��`�(cPRa���-|�% B5 (�&鈗�Ĝ����Vؤ��°kW~;���{��������b3LR�]m�~�d�kq>-�oP0nԜS��G��(���w�Jc�Q]Sz_������eIDɞ|�Ŷau"�p�	�כ�l~K<nmI�D6\�f����&
~�J�����v/I kڐ��c1w|�y����4�7(Ǭ�o'BS�����C������%r-�(�|���!e�s������ȓ���U�� � �2I�IҶ�+;G2x��۔��3���|����"�W�n�o?��2i�O�@�0t�ŉ����gF�.}�~S��� \�wjh�oq����(a������v���n��=!m���:Sł灺��0-&sD�� -E�Q�itA�wRdr�z��{�?�=-��5�LuE�b�6!�L��1J�r��m ��R_f��o�J��E���	8��\4)�j�͚+c����!�E��{:S�|�l���y�nn�&Nt�x`|Uc����?�I��@S����FJj(-���AdG�>,�[
<5�i��=ܥ��Tv`-�p<Չ��U��j ��z��3�))X� E�����צ�؄2���L��ZR�\����nx_���}�d���������ҝ��"4AV>�H��MH��4���%$��9O/M�����Z��"�1u7>t9vf+:To+�O�+����`�c�ni�V���m�S�=��Ir��fCP���R�y��&�fi5���]"':&�K���s�gPed�`������x6�RG����=K�Q>V�h�
&6�#Ov���&K��+����1��#�%��g��}"q�8w<����i@I��>KϾj5�qK{�޿2���u�H�ɯ%י��W"���FY����h~���焎!DV�9��v�1'���:d��C����Rk��&���YZ��A�)���S��ER���X��� ��&���G���f�l$:�o�<��>��ƺ�,%�e
�F� ��+e�Ի5U��V������}�V�WX���!� &��H!�'d��0^G���~n��|7*�-��EA�_�]fX���_�D�aD��	Z�>�!���\�b�����,�9-0��рN"�I�2�rZ�9���v��M3݁�7�2���P��4 ��#�=�FR��(��Y�H��^Nu�(iфp�]����2)y{m����s��b�����O���'���q�b���p����˒��㐎��������e@��\�d�IV�#4��r�����\�vh��P��L㸛e��$Sxbh9�f/��W��Z��P<Q�;��,(/ZG��P���N�;�����7~�}�6<�#"r�L��O�G	��c���֏���H[#��s�O:���m��]�Y�s���.x_ǧ
w�Ap o,��r��!���/�'����G�S��X�H��^��*�Wy̅�e�B �K\M�H�[n�k�F�0�e �<��=���	�W�3��0`��X��3���R�E���>���=�Ϥ�Ј�fXW�����Eq$X!�&�֎{kqz�/��P5_�DL]�d ��<�:c�v�Ι^�W�a��l�ó2�!����kI˱,ZB��z�kP������!I�쳱�~�4/5��=�.����L�\�}�ʔ��L�IgJ]�.�pZ��D���Y���#dW?��n
m>�7k�����cN�c���I�킛9	�D[�JW�\3�����ՠ;SM�2$�� �7Y�"!x����	�/J��f�|��Z�s&�3;�
�)�$��	fA���.���C�$��e'����Fd�T�>�[׈��  E���>�)-�Vs)�]��/�a��>yzn���r�;�CS�!��*�O�o���:��x�}��À	7>��p6�j�Er1�����N��[�%)��"{Ŝ ����>y2 >�g�G�:��Q[����	���d��b�1i@���5!�����{�_q��iwS�yN;d�ۧI����#�~$m�m���b'�-J�)�{@���Lizh��Y�r_�e���+���KP��[F,�'�0^?�Gk�䦼�H�b5�,�|ڧ�"ԐP��'��9�O�����[I��h�){���X����}��faT�;ܳM�G����!�Nx<�(/]���ȕ.���m�8 h��;;|�JW�b�w�5�K)��s�?�}0G}멼�ϨMhc{�a���	`����//;��圅}ҕd��;Gx��$A'�ْ�2�RZ�?��u��媎����`�m�৺玮zͨ��$agP�X܂nV]�+�S4�|W�قr�Xx���ᶂ�g@0͇�]a�b����,�P�)c�� DeŜT#�{�˵�ߢ�,��������]�݋�p8l0����]�P��zQEϦ,�T�r	qGX"�¿w�.�`��������>�U�pb-+X��0��*��xu�j�S#PUu�V��$3p�Q��y����OA��u+<���jԥE`�.0]K ��B�P��_�[	��{�h��{�����`�|�A(�oTզ���[He:z~�֮0M�,x}�LQ�lVШ�VH��ey/���a���N�#٢���X���H:g���U���Zhx���:p�w���EU���cj�T���H f���#�C)ߗaY���RM ��=d��B�ͱQ�Į���V�z;nڒl{�x֠���q�M"������lϵ��cU����{��-z��ə���4��^���ȕ���K��:��� ���9���yX�w�>(�ga ��7p\Нș.�ikk~8�ȋ@k�J�
��ӡ2�$v<.��K�";k �-�U�s��F0&P�Q���KY3��E�C�u���G���Y��6&��>�\��y7��N��L�|��-T�Ս��;R�x4���<"�/�F�'v ��I���O�P�g#�����mc�m�����RF�U�d\�E��qC����+�A���s�bPAѣ�( �2��@�}�As(��T��fs�l�f�}$�,�6-�{|�j1��O��T6�������1ku�$"��@�!H.�<����Z���`КRT��[�H��dɚǥC6��.�R A{����T�3H�>�iS^��a�n?k�ѥq�@�o��U]&k7d���V�P����VV�u#���5�ӥF|�ng��҆�X�bGX(]�O@QXI���K����n^�D ���͆)�K�R��̌�th�o$�܈�62���̆fG!����[����<�f�rH$b�W�j�H�W�s��Z�r� �U+�x��8�웆�}��b��Z�ph6%� �1�}zqm�_֧�%��pnoU%S ��K�w�Y8�杞�ыa��U���E"@/�%~{F@a[&�7���x?9�`��B˄�T!l���:�ͦ����i<��b��'-St��b5Zrt��dC@��Q����pﾶ�*5ן�Y�������2>P��i\1�VRZ�zc�����)���P���-��fQ���2�_�@J����]C��pDy4�G��f2�U��&�6�l�������Bl�T_+�m�9.�D������gՓ�l�
�[�>n�[y�`�4��Y����b�΃�� 8M���s���k�b⛻[����fv�9�lQ3P['�R:�z�д�7j'I�>V:�;�����%{j;G�Y���k2M��]
��_p������@�K����S�p���iY��q�.��������`����Y��&B�ɹ���0i��� ������6���qUz�7;>{�!V���I�lB��R{�L��#g�:�R[�f]���H�a��jN��j�yʢ�A�Uj�ӫT�<._L7��%��k�˨4�"g�^G�������&��c�jK{�K���Q��1��c+��i�����eM_<��Ғ�!v�z�����ڵn��e�N.��j5�$I\�el�����"e�=|���^.��k��r��6=�x�������}�<�>�}���sI���tp?���k�C!���(*�)<<>�D�]4v�	�
�zr;����G���}6ɼLW*�5"yʽ+�-ӑ7F���\�@��=�ǎ�J(��!�.��w� �tg�w��Z^Uȡ�Y�+����'�{����Om� n�;١��bZ!Ҹ%э��y��3N,eZ�s�|�& ��jQ�$U���}�[yL�	�Sx��]���=�aS�K@0�I�k⑋Q Z�U�|#�0��2ή�{�ڀg�l ��T�5߄�!a�"���4��l�|�l}E1�7dCp��r�Yد��7���Νcs̽}G�oB����ځ��y��MHu݀;I�}Y[0�U��=�n��\Qd�S���|ӥZ1�v�1(���C�k~��\�s{茝�������zj^���k��A��b���GxcO�������K���.�|�2�`�Od��U�����D�w�x�C�wyZ�]���g��Ή�_�:�y���m[���%m,Z���-Q��bj��F.�'2��X	
�n���.?��2/d*h���3HA|F�ѧRN-�v����x/�哏�V�����N=�c�բ�!���f⦇���	0|������n����K�e���n�e�t�/i�9�����B�8YHi�p$�o�+��Y@DB���"����І��R"m�j4�h�(`F?i�S5��Y����q�Irb�8LP�JX�v�;e&XջF!�B��HE�Vf%tb���i�v{�7�_����Z/�@�!ݕ4��q!J����$;��j� '�F4OO{�?�3<l5������x�>,�Ib�v:���Kf�+@�F4%�����υ�����*o)�F�k�W��QZ���q׉� x*�q��u�W�i�@�d�ah��Kog-������e�|�s~㜧��ůR��h�����6x�ҋ�����{_}�o��'�^8B��@W�Q�Z�_O�<�n⪺Qp
�������%�,A�b?��gӺrw�@2%�8�}�Z?I��ݢQ�WFK�$��k6�T��ڹඎҾ��Ņ�&����c�&,Cmj�S�1oS�M�6�7Ѹ��ء�;�Q�hr�����~����<�d���b��LH��q�������݊�+�0 �p�M�Jn�*p���_����_
z�ˌ�u}�t��Xb��:i�cg�'��S��=N!�9x����;)K��$,=��2S��S4�=�xe�zf-��	i���ߕr���$�z�m���%)����*�� &���ZE�c�x���x�qj2��rRQ��i�y���2A��jxD��G�l��ꠜy�U� fSx��Q�^1a0��9�ӳ�
˷��H\����uM~n��X�������[�p�����6�DG���S� [.��Uu|4���:�ߺg�������L��eiE@���=E��#yE�M)�z��g���*V��w}q���5y�G���\���Q���a�r�Jl�ܷ��H��2�BTQI��\.���]4-�O�/��O�}����%�f�!Խ$L�̛/�AА�n���F���.�uUg�<Z<P��)Z��y���F|)�:�B�������l�A�A�Y}��u��!_`�	����,&,19��@j�h�	q��4���*��9}ʻ�����r�(w�f�S燃�5��_�~���>Y�{�щY��I-�l��tv�" ���#u�r��������3!��D.��&H��Ͳ��W���,�M͝Cύ�4iP)�Y�ڿ��6�3_ћKQ�i8{�ډ��#"ŪV1���(+G��m�*݂6�bq���C��S��W��Xϛ)E@�FU(��ۣ���}J����J�}}c	ƨ�2<��#㷹"�z��8؂y���;��etn� ����� H����g5�[*J�z=��P1��>�W[̈́D��<�zY=�d���9a�\��T崦n�7#D��9�Ю�Cm`�����O[bş���%�W���{{j/GC��5�#� �Ye����Z�zDU�D�+���R��`���8V~A��#�<#���b��3q�]l	|Y�g�v�>�Q�]��]���.����S������IR2RcA���nԇ�[N������A"�>���qz�!���n�����XXY��9��7�e�I��}���nwʐ�f�d�q�P+P ��r7*�`���l��D��x�4�p�3��8�v��p�"��W��i\�]|�	���:��C"$8��9�ï �O�=L�@�ٵ�)z+� <q3鲥׎���YS>;f0�F��c)g*�g��(#��a�}){�4�������o
f+e�c��afţ�#_]���2����9tp�3!y!����h�|��]zL��BJl:W���Ǹ9�^�I�t�Ȟ}��\��y!�N���ƚS( �h+���wR'"��|�qi�D�r�4A�����u�)�_��qoYڌ����Fe�2.����M�zˬ�J�+�a�L !N�}��O��fA[m��<��R>���ˆ�?�s�B��8��:���&�M^��xh��ŧ/'+���z���|J� �K�h��ւ��&(��F�]�*�PGf!~��B�M��OT�����s��S��B��9Lv�%��c%t�-ߙ��ǚ!&��YEL\A>�!�w\v�0=.:���X����vB~��i��XV�,dİ�N�p��}�t������[�U�rD�g����*�T��vq�B�����∹>�],���#��\H��lx��<��$��=���.�S�vJ�x����#zE7�4�uV}�nH�8��@�ӑ��[1���� ���C�?�������E?)<Y��y�b�S�=�
Z�]ߒ��
�7���J��x�'@n�`��JA{`��I��W�|�R��п��e���L-1�9����D�3�Ƃ�lA�v4����Sյ����P4B�`>�Dڬ�BL�z0�-��áSk��\��Oo\�`G�4�<؏BtЏ;ݠ��S�E�c�!*���&%}%�����<Lǒ�H�OL�Qu3z�hʑce��fM8 P:5+���Fk]yґw����P�}]�~�$���'�2�'/#���v�,��fT���������7�����ݶ|�[�W��X��ȢA���w<rR�K9�� �(v�f�c?z��I|�~ZA�xX�W�;��j�8���<�N���^먚4�V�^GV{��=2��+��3*ʃ$O�N�%ǎ2���v9_�(�����mK��_��I���`�L�$�X5@X�>�����E�lc�;P�6�T��J:�zw� �rw�B�EY�30{��,1�P�igs�����~9���kG]!ז��ϸ�MIV21\�:}�X�Fh׈� Ma��l]bN�Yl�<�c,��"��\F����CN;6jy�|WR/p�=� �Mjhf��Y(��B���c0��4�jd�B�jm!�Pd�l�z���[�8���>A2)���޶��[2(��2�qђh��g,lY�8'�K��&���|�MQ�,�	�GzF�봅8���E��-l���a0�.�������-*�l��<���u(����9:sJ� ��|���>�L�O߲O} �^��� �9���`��+�R�/[��d9�1KDcK��o�+׳8.l�
#�.��jT�L�����Vj��ꢴ��b��b�^��� �,Y���Vy�\�0��MŨ�A:5%)z��d�}�S�)�-I�*����x�<��J��)қ*ZHY�ln�/�@L*�N~å�٠��y(>���;�O�I��E�-br�;L�L�]�H�qrJgQN���8̂�7s���t!���	�ڎB=���Eo�8��܇CY�g�a� �qk�d [M}5����P�Q�����l�\�
�=�D}�+���T�2O�h!�3�+&��֮�*�'�G
�b@CE���1�;�	�	+k�+��`<,����W����Q<W����!Pb��W�̈+q���S��o CД(O��m���.w��� D�xL͋8Gf��3��\�cbj	N���Z���}�T�{��*���v�zl=<eԙ$O:0�#pN����P,K@=����A3n�R�$�Y��M�T,r����ꩭ���)��Id���3�~�����*Բk�2x�����qߏ��?�)�Yg�6�'|n�l{���x����m��|��*���)���!l��w�:3k�����#�u90U������Ƣ8y���|Փw�x���y��Sh�:3��� ��mdh�{�X�C�'=�ǱI�{%Q�~Z� Ot3oR�3��C���2
-��0�^x2k��Ր����@�8�����S2�(g��}�ܪ�%�XdSP�4�۝n���������Yc�]�����$�4�B60p�o�;��-	ݪ���(V��s,��j�ƛ|���.�;SQ��~o+�Q�%p#��ͪ��H�t*���]M�9�kv���_�*;�X)8@�=�>i��T�? ���R�` NS6���cY�0���/�2J�����>^�v</
'gj����V��w&� ..��Fդ���;�ˠ�0UO� ��e��J�9��6�n">^*Q�f�P^����[)�[�%�g�����&��y��x�q �����f��_s�@YT�sy�v��;7w�!%T�q;���?�����E|9|�8_'U��9\Vɇ��W|_�M
�PN���2�I�b|U4q�:�,�1�_	��+�#��L��_B��"7�o��L��V����қ���<l���E�*Ͻ��G=�7�˫/j쯖%�T�x����I���쌈��WH��kI�2A���c~C��`k��;���c��� �&
���kJ���AD_(q�/x��(���מ�Z�1�����`dv7XmC�ZK�߄ܖ ��<�/�k��d8>
X�����Y*���z#\��!�x4V�&.�������N�|f������汭GR@}�Z����n"A�Rg�~���cm��&' Y9���� `���vV�o��p7�MP��e�t˴hB��1b�Z9�%K�Ak�~%Ʈh�t�_5I����Y�?d���#,o�9[�|­���@b����f�p� �A*�1I� oM�QhV�����K���Fb�r��Uu�����]N�^�	B�+��a5�D�kC�Ў�I����E|�CJr��K�j8���V�����	�g�A�K��]���p�׃�>њ&��L
<�4�6�k����&���]ed#���h9���t)M��O����H��n�[M ^�0��=��3�.g��K�$������2��r���	��{��d<6�ʤcc]4�b��e.ϝ^)&8��9�a��S8�;UIzQ����q`���fQA�fv֢�,˫�쥝��6�,�G�/�G:��'�*�P;�K��>��>��w�ܞ�&6�<�	%�=&�1��#E��
���2ZF�%�O귑�n���'�&����e����$a��*�����F
��/P���A;�2%qq�u;�j�ь�fc|K�z���jq�	:�c��{5X��x4��J��w@7&����S�f�M���R�m]=am�P(�bǽ)��ԘŞ�������LQ��P�����}<v��WU�%�$��h|h���n�T���R�J���"
=�?8H1il>^�TC����$�f�cG�0�*^�5-*�WL��sh����ONYI�r� M��
�B���=cٞ+��U�H�7o�*a�����Ŝ�o�7dsV���5�[�����q��u�ڌ�`J���΂P)�&���i��~��9S��rk@${C��%Ab���*��>ߩ�W�to��<λ�d85��V/�pPNq�%o�s�c��Y����w�OJ��}�V$��d��%mc��X�YzQ��͑�̻� ��s-�y�n�N���ݺnm�F�!�w��Z+�2x
/������7�ֱ�-&x�BA�}�p^0�Vv-S�Ok�����g�	V�AW:P\���Hɋ��ki�;
��� m�&bT�딸��]W����j�]I��r=S7���eo��v����v�rp�/�|]�w'��N�&�+��}�%�Jb� ���I!�T��Yh�0y/e��D����Y`D�T���Ž��.P�>�-����H/�� ������1$��vU[=f���9+�������WM^ű���9��1��-�ܛ�)��G�=_TuCӴ��g�o|���>�	y�BPo�e�>	]u���}g�ܫ�B;� Ɣ۰��?L��{f��@�k@Ae��̥n��@�3z#5�yy�w�9�J��'}l�"�8O��q��	9ȝJ�͘o��A�Ѵ*/EsC� 7:�V�Lޝ��oH������|}�ݵ{��z�);!r���p�`d͞@��;o]R��Q�׊�zAL�\�+���xC^���0�mR��8�^,�	�Q	���t�G	��h�����9E��	��_�x�ԅ�R���R^џ.�h^fR�5(#'�ZIg!u�{�8'�G���=.m�z���I�I�������f;L��� ��"Pd.��C`��u���z��b���<��|���ay��!��H3���(�X�b�8�O^���c"�dCv[�W R�4����T��̎ງ�i{���e��򁃱.̄v�|p��Md�4���[p��ў���소~��5�4f��s��o2�Pp yT�=��k�.�!u���@�S3et6������w���Ju;�5�l<o�w`�U-�-�{
k������+ab�)=��S�o"9�8��w�U-�Y]�� !��}�u22Ǳc��:�y0�)X΢��S��9�K6�/�f��}�J�۞�HWnW�}�FQ���F��M��1e�ZR;�\��4-$g�5s�7�h�_�D�C���C�HҢ�,���=��4#�?^'0s��!�?],.5P���W�����SI"��Zx��R ��yD>[Z�e��!x�f���$��W���{h7}�����X��{���vWHlR�|
�7w�s�l�Q��<:��Rwo�b�?�6~�ˤ��<���R�\�Ђ���,z�}A��'�$�[�i+Φ�n~fK�9�Q~����[չ��%��~Cu���P����~.,���NR��-�j@�;3'4)��R�v	��3�}�I�GK��
r�&���,{�Ԁ��dI	w��(ȱs�wH����	0Z
��p�z=�� �b����(!���뽩K���h�j��m�U 𨺳3}�+g'b�@���깏�%�����?s�NX���.�Ȕ��x� �W�s�`�~�%�=xHo���Pެ��=����bT�Y�����e�W0�|ӽ��n��m�TyU�?�b�z��]�N�]��M����ɲ�>vx�Dρ"���9���T�G�dg��Ywg?�2�ֿ��M���?*Q7�3��S�W���I�![-�� k�`����Э���?]\ܐ������i+��!L�����pj�@�W/��%�ʎ� �O�))���ti%�}�\��[�&/Q�D$�j�ů������E�;ǱdBF�M��E��e뀟[��k1k��5��^����T��v�|;���7�^/��<ᓠ����@�����L��^>#i�0�D5����y�v��rP�{<g��G�КvZ��vL]�&��G����xj����$��){�Aá��΀QC#��M��e{���(!����Б�� ��'���-��a��d�UETs�Dz���L���u�����35%��ɬv�ǰ��^⺩�A$���) �r����>�S���t�����7J��0j"[M#�6˝���L�t^�T�����k�t�h��H�;r�a;D���)p?`�wy�O�0�X&$�8����I�m�hr��D���������W�~�I�
R�v�4+��my�϶읿WoT׼���+��̥���N,c#i�%Q�߳�47'������%���`��-����n�q5��>�	�xc��>f��t���E+�A�,w�L;�A�\Z��5@٥��MǍ��}��k�J�L�a,4���=h�\��Аd���*��#�%ԓ��HҔ:�)k���a��?8ټm--����M	
b�j6��~o8]��he��9lz����	��ac�jx]�K����W�^�H���pA4@T\=��h�����J���
ʾ�vۄ�cG����1P�uT�g�@�`�fcZ��:M���}秿p�B�4���j]	�c�i�Z: �WEk��I���(#�
=���a"vAqB��QxW��#8sŦ�|1�vð� &Rc�����=7õî���6!{��;'�-Oj|Q����x�؏�n�S�_�+�-�u�%�8��Λ��G�܎$�����=���jp��׆�)T8�@m����2�u�M���z����~�������o�B,`�F��WP��1�MW��α��|�6�Fy�o�t��9.N��}t2�xG�Q�ֆ�x�;D|��14V)mK��^��Rw5�[c�7iF����8���o
oy����_rlT����Q��(7%��lbYk:N<��S�]�v�B\�<��q�7�$.:z��(]E�h\�j�Ȗ*k�
@�;��J�x������aN��Fh|���k���m�>`� �{w�
$��Q���?����m~N:fc� �ᮁ�M�	!�J'�0��@M~��)�����s�,��ӽz��1\d�$�/�
]���RM!X3�,5�sQ.����"��T>/��j���$��pS�Xdf�?v������:�6�hw��.@����ei�dM)3t��Mt�
��u8�� �;ϽY�X��:�ೞ~?&��8K�IB$`Xz&^T`�����}���l5���[�ov�߳-�0w���V�y^nj�C���0h �+� 	��weY]�m���#�F9�LHۍ�'l�+ZX-Ng��K>�u���P�!8��
���� �+��"p��
�B3{�s��ނ��Ѷ��+�s|W}�xX���7�6ݎ!��U��XD[�`)đL'��I���{W���˔�VF�� ��O�����]�XaQ�:ϴM���D�pO�l��q�R�;y��R��Q��W!�R�W���Ѐ�l���[��0��i����"���2�Y�3>:�������)�n���>?1~��Į�'�Y�K)|�/~�.%��L ��Bʧq+�L;�F�-@E�$�>�Y)����l\݀0eq��7��ll7�pc�灚ٌ��[��D!���@�u�l�D|��
�31v�l-eRN���w������$/h�:˽�\)��X���+;��ծ��κ>�+`��h�oD�
�̍��U���xi�N�S�"[��+VҦCx����ȣ�����$u��B��t��k!~��	���a��6���Z�>=��~��Q�&Ȭ%|Z�/O��q�Oo���	ID��Y��$¢����A�L
�T�} {|9� j3:��*���Xw�9rY��R��B4���y��9�prq1b�ϯeHw7M=!�A��B6�F�_(��)�[R�x�8O�M���Ib�/�/!�=/��v����m�81�2黄m�psI�S7�)7@�"�*U܃uA�ʩ..������v2�8&|��\�7��)�"�x���_���������G�9�9_s�q����7�$�d�NR�d_S�XN�e����nC ]��sq��0�g��i(5E�_[�ԵA��7�#:�����"ڭo7�����S���p�uQ\����a`�I)�t����qn߇Б�Ē4�����`M� Uc'׉ߣ�N쥃-=���s� �`�� ��Ʊ��֦�.�(_�{$+���Y�v�P��7+tg!�8ҿ�i�`�a2]_�PI�ov P�ϭ3���}����;EBk�����%��FPMj��E�ߘ��Z�
���<�.U$iG���:U4ny�c?��i���2'4�5�	,�O�饷�RW�U'���.;OTS.d�V˝��u��w��>�����.�}uаA�!����_Y��K?4���a�ϗ�*�x�OL�.n��C�2��1h���:;��Ҡі���;���6*R�!�Ci��5�aZ�ML���}3B�(f[�:��͉����7�ܮ���]�����K��謢#�=G������̟'8A�� 膽�� zx�����W�a���n��GAe�i͈�40��%>�-�+,�..<���*��N����)����7�V/�69�Yg-�z6No�ws%Y�Ѕ�(��	��\�1�)�v�U��T{O��n/+,���]�
�0�5G�"L�%����
���>��.�k	�C��� ��đ��/�����.gE�g��H�'�N���H`��?K?��l[09��^0�[���@-Q�%h���+[F�.�*t��s^�y6>��)?�Z�7����%�)����WƘ �J���Sn���z3�!7N�����EXA��3@��Y�RO�t3bb����y3ċ��G�ק��A9��gW#���B��<P�ݖ�ia�ӏ�� �4b#/@�摂-��/m���Z��m����pyT���^��caL�1���O���a�s'R�g>�i�=z�iJ��Q8$�����|����њ�ƛ]]�}�������Bo?�UU�}�j�Ry�B颜��.i� �z�kW��u3x��!-��4G��kv��]�ȯ�-47
A�<h���{tB!S;clHkP�v~�'�޿A��៣�E;��t�ξ֔������ď�Cٓ����4j��!DQ���F�k~��S�}���#���	�u�n�l��-f��Bm�zNHJ2�U��̧+#	���W]P�j55!~�usY�2��w?3Pt�n�F�U�[KѤ�D��U{�]�h
��)^�����\pe�d���V���_s�Cᮍ�e^迠��[��T�j����}��Yu���3xP �
ϰv�v]�X#�ڼ��o[B��֑~�g����t�{�`mC,��}"�n���nFF~�^������)�IFB�۲\�d��U��9�Q��^4ۜ�b�Vf��5�d�iyI��'a6��� �i3;7~�L��L;�M�a��K�oP����M�SM�ˉҳ�����]�Y6�P�����<G1��u�5��M�o[g�!�y����ǋ�`_r	u!@��>�,��ޟ�E5�VtaѮ١�I�5�}�/���y�"3^�}��OHqt��:I�"e�vX�|akk��z�����	ȑb���M�;�!F���C:��������4�M��Y�ßZ��A���H%�a� 19z�ɩf���X]�ׇ��iM��j��zm_ �i���S�m�d�NdÅ���',1����T�{Z��A��:u���5���B�����%���/�a��I�H�} �H�Z~'t��cX�>�����v�}�\\��S���M�`�D�HGI�YqJF�h`�,��@� G��{�Q����
 ��=��E�&����$s���%�>��|b�t�.)��	Ç�9�B�Ϥ����w�_��9Ic�������x Ӯ��ّ��?���S����~j�?���)�G���5�^Zx���	?�*oՐ�����僩Hvώ�'L=�F��I�f�u�Bb��(!&C&�z���W�w������F7���}�7C'��34r��l�K7WU���V]xP�����'{-�/jS=`�bj��E�{���p��e?U*}�`h�`��@�NZTv��QQ�Z
��k%���~B��q�XIs\�'u@[a�-M1EE�#��ɡk}�Ř�͈��o���dT�A��=����Brt�>ĭX��ՋA������*�/����6�F�ox	�H����aD0Gr[1{8��m�	ίJl�LO�ۇ�*�Q���@�)�$H��d�Ňu\Ԃ~�fm(�Y㼒95��<�*�5P��B�,7έ�;c\Qn�َ�?i��8_�h�g�ߞ��ۨ �:2� MsV6r:����菁�ϲ��'�hn�z���8�����������Oc+r{V	�s�#���ĥ�i����0���LI�EK�t�^�S����`꺝��QA�H�wW��#��Z�1?ƎZ�RޚX㻁����4%�*�7�Q�̩�� g�ra������`���J��²���>]� U�k<l��n@n椞����� ��y�
�v�Q���j���i�"1g�ǵz��?�� <����|���%N��Q+��α%O�u@H�hW��$���^6�~E�}]��M����/���S�h�����zd|��� �
�Y����z������F!=N�N���xs�\x�}|���O�ꈴ0V�<Sm�T��C�����`��
���m�9��q&;���8��#��4S0SV��*��կ0�R�z����8����XŖP+�Z�HEU�N����f[��?��G�ȾT�Q	�c"X�Q��V�f5� #=�Mn,?��HdU��ҔnT�Nk�%�$/�Wz,��Zʙ�D�	d\V3��`?�Uv-k*Wd���4�u?�6����Z��5D/�n�����$�;�G8tm�
�Cn��W|/���[D�0?q��9�M�2J�uk8������������k���9�{+�(g�%���Y#��ְ�w �a[Ur*��n"��j@Q���f &����?�#��Kq�Z���,v����.��4�$A�a��P��V�^���n�W� p�6Q���0<Cp4�N2�.^���?��y���H;�I�ݶiA�8M��-�����+�a��V2�5[����F�{47�~ۚ)R��e�HC�l�{�).��{��V�`S����錾�ޱO��]���P3��r�h}�n��N�����Z�-�q��?ӷ�����O5,�2"ҍ������;�����_FJfU���>�ص��f������tj5O�HO���f��w������)a��'�f���7��E���"�=vw���/o�
i#��9G���&���B����SC=+�	w�%[Q�鍿��B��Y70g�Nlպ}:��"#�0-<�b��^���=ա����/�r�4߭�Y�B4)
��F/�~K�nuzӪ��֓�Y�y��UP�f�}��ǭ��c9�
���诔���DǾ�-�q*D+4T�E����W���|(��������]��uS�Ѯ=��Ρ��������\#��R�����9ӛ��z��fG��y[��uGL9@
�m}
E�&��ˏ��f.<�O��	&~tA�X���^T���ryź��H��#�}05���RM[��B���	Qr������1͗>���wК�;c�\o��n�� ,������"u���^��ŷ=����ۜ6Pt��d�ǈ���/�Z�ƛ�1_Yj��Y�{1�ϡ��_~h���ȸ�#5ɥ�0��@P�c�UL��#E�!���I����ǥ�B������	�^�<�^
y���D��R���/	����{����>D;�D�3��[бr?IuApK�nc�%�e�YF\�څ�ȡ��
���`���̠NBuax��tա�m�ѼaWd��( '�`�����R����8���'�'E���D��;*���Y�h-���Q�b�v*�uv#p1��!#9�ǧ��M�]*E>۬Y��呟'�&q�^��R�?��1�aQ@���4e�k�g�C���?�p�\7�S6�#��.�^�,I)JqQ���ɨ�XO�h��R���t�b֫}���x�k&�F���	+e�<LmV$�`2�z��ӄ&x�� �3aL����90G8@⹿��~��1��x\ĵ���N�	Lk�CF�=��#<իX��,���n�M�vIﶄ�q�}���� ��J��6�fĆ:V@����"��c�X�&;����{�V9t};������X���kH��[ymXP�@�;fNl��?���te��_9̢�k���o���	z֘H�,ee��o���ou	��7�"H�U�*e
A<u�6Rӌ��N[��u��Fj�D�Q/��C�[�-��L��4�����0���#G[Ա�Q�Z�<|�uО�<�x�M��F���+6��i)h㫣���-h~Wxy�S���B��A���Rkx�[��oWC�ge=��:=��	�)��~�}���&��&�D��t������49,H�4�nJs��1�-��'�e=�-��_o�W"������XY��e�-���irC��JN��ݞY���s=��vx
<��J�X�d�:nA
���pּV �T[� �7���HJl�Y|OYN��&d������t<�����uF��-�U5��D��_�y�X��<
q��z˼���͠�ogq�;b��s!��~�n� 3��$fΌ���R�%-z-G��]�DI3�������2�d�9C���_ ��79뻺h�GO�X5n7�}���>�
�6)"0Њ� ��n�I1����V8��ڋ}(��'�|�OS)����fྗ��61j�u��('c�9��ˏr������5	�+{�yr!<
~8�9���g~@o�֭���U΅���w����{�o\����g��u����J۞��Lh]rb�Nf�ڵ(�h�eŹ%�#-��0�k��4��Jm�t��~��A)�U	0%�w�4�U-B%�IF&]�n�9�|��]�Ϻ&?KKLI>+�V5!�����gq�&Z���5�I�d�JM��ё-�$���۶x�2�.l
"Ļ�!���j:D, ��zO"���9������9O�(Bk�(�4r?�b4��)q�S6�T�����X��4oԌ����x[�p�����ky��g������t�c!���@xpf��̚r�;T�g�w��^?�@�%]���+zꓻ�l+�ȾN<I}�U[�&��y�~�cS��#b(?�>Q��:r�=>��������
�i_	1i۾�|�M(D�����뾠G�3ŭ���V��Q��s#���]�������#�B~�Q�ee:�U�ִ��W�Lķ����t�mX��my�^T�T`kџش���<&���p���6-&.��%��BC�@�����DL����>��MX!�5�*]~�o0�KF�H�<�X��fM��UĐ\18�h
�]��LÂm?u�(��z����b�*��ÇhD��<8!FI��d儱�O���u�b��3l��s��V;���Z�L�;�,O4`���H�����|��^cͳ���i8s�V�Sʚ�o�9GN+�>*N��Zo����'���`9.���TM@��rJ����Li�~RR1@����1���v% ���7�K�F�$�F�[\oO`��%��O���-��Et)-e�`J���@�ia��;��������Y�i1ܦ�ԵB�?��0�J���6���Ün�Pю��6� /l��л.�H�G;8,��v��ȫ4��Vk�l�'U2'P���:���	� ɇ��ɸ�Ul�_���	rqx��r����[��"z�5�Tw'�:Iĩ<'��@g�5p�]n3v��[̇R+�ϨIvG����&3+Ij��b*{O�r��g�;.v'7~��e\c1>���E �i��ruϳp �-��:��-���I:��Ǟ�0D����������O�FAaU�E!#Q�F�<s����4�h9��GjU�i2�X�rU�wI��d�|�g{�bg��'�A
���Q�\����ݲ���.�����ໂ	�Aը��J����!����������m��}�&��郠c��:a�Y�����Y�ze.����-����������?�w��G�X�_�MoF��R	iyr����:���(�~�����x�G��N/�!�9-&j�����%?�h�l��dYo��bb<!���b|�JT��Ӧ�0Y���J��>�jHZ�&K�\��D��Z,H������bp]��ÞJ�[��O�",M ���A�NV��Q�e;��ꍔ⹐�鰮8�'�,f���ZɆ�B
��B'\ԛl�f��!,�m����SDg��0`��M7��`N�u�(*Z�m��sF�B��N�F�w�Soaٯ�Wߣ<�pK�������:{�`�h��X��o����N�T{�,�TA����+���yޘ�WY�y>5�����[��H= ��Ăb�|o����Z2D�|1/}�����EQ���)Y��#��X�+RX�����f��Mqֱ��
n&�Ӛ[��"�������`w�_�ҝY��K|�tw��rv˭�p?>:���[I4����SpN]�Z F��҆��2Vu��s/>�ʅ�{�]�ͰJ�*�1^�E����ɽ��~M�S���R�	±j��ã>hѓ�²��n��D=���fΦ\���b�� ���ul����0>y��Ic�˭�� ���8�K�~C�X��F��	O.�)+�9�閡d=a_�5b��TUVa�oJ��|�I�?��|j}s"���������Lde#�vB�E��5=�A �痪�&T�)\{��5?�C���k�Ӥ?��u5l�3V�}�T��\O���2�{5�>lY���bH���0ǨXl��y�:����f�=�������OAid��cǇ�����Wr�k2�VùSN;��!UJM�{`#�
���$�CPiᆕ]��&��Y}�>hɣK����E���ߔp��Qͳ҅��dk�H�k���ٮv�j{m�I��$xOS��XIQd��yg$|o�>%hA��� ��F�ؗ���C��)aK9���W�;)�Om9,�����)T3p�/v����͗ߨP�7}��������{Tj����- ������ܻ�N7Pʾ���9�4�O�<�U���ܙ��u�,�Կ:'L��	O�ޣ���q#���_�$I���4�c��hH�S�3m�X�������c}��
��R�R��7	��7�$\L7\����c0>�T����δds�T �;\��u@,���,�I�Tm\`^�U�M�\Y֊��z����E�'^��ظ4P�X{�m/�ɼQճ��5�9�2�r[[�;PfHGm�4?Y�!�����{���?���sP���3Opa��Ψ��׆�UD�iqG.EI2" 9�f�(���\�/�ŏ����d���8C���}ƫt�"sԐ%�B��澑u�^�ʨ�{��ġg�!�ᵞ��y������Kh���n��Y�(�? ��Kv;��E ���
+}|fA�����c�
Vv\�(�:������� -�W�0xZ�,��+X#��W%:�~�0q!G��n�#�׀\s��.�4�L��4��o�.ז|�5?HJ!{X�h�h���-����L�R�<L��������6Y���4)��8ݱ�E��&���,e �k�8z����a�Q}!=��,$����%��Xu��J�T���r;)m�02��/�~��7���M���g������yT��T�L� ��T�^�t���ր��!�8����t��?d^XS0�_��G�_�i=mH�]��M8|7%�S�J
�i�S֞�>��A����\�W�60�*�<�[��$K��qss�(��a1v�T(��s����|�d����2�d�A~�x����7�,v�F����p��D
�$$�3�������vm��q�����jB�U��`������z�����4�Wg\�w״�{	�\��~=;dm_��w˱io��ahD���P���k�m�j�'��"��ӴP�c_~['���JP���O]�snX�l0���!8�Fn�"r�!�
,���S���/��bu�~�g�����py��S�͞5㜤8$ ��,��2�f�%�H�	�G0���BR6H%Sk�!�uq�ǯ����U��������&|����ª ޥM��{��]�&+�+��Ҫ�:Ĥn��0'�#�T:�;Ed�R|����o	�x��D4�����OS9����_��&����V�h�N홄:fN,[�L�R�D��>	�@�u��]t7`w��^lM��_.>~���Z0��ّ'��q��t��ꙟ��T�؇�4'��A�j];�ۣ�-Z5��e��3�IL�&a.Q�>��Q�.I����Ҫo�3�P㒶YK�����)?�n�U��My@�OR��f�d��T���	`̸�G4�H��N���nI��^��Jɭo|b�_X��XC8Oi����zΎ*R
�g"����v���M�(�%)a����l4v�j���=�Z#Jh��d�b���C��ns��S���r��t���*�;����x��'"T�J����5Ӥ���M��� d�I"�&�� ��U��{ٿа�����e?�"���C�4up��C�aׯ'3Pѿdkjԩ�+��������<|9d���_�!eF�� ��+�L���%wk��@�i������:���q�f��u/'��Β�}:M��r�!���������ߪ.���
��gF:��\R݀��{�d��Z��C*e���sFЮ��rR�
ł�$x��)گp�C�b!��,��?eQW���L6X�m(�S=	MJ�^7|^Q��W��.���~���	�'8�<�w*�$����-8���DH/�8���N�d.'���~qFn)ng�
=p��������8�������ن�d�;���l��v��A� �*0?�2����^��Q�hu�	�nҙa��F�V;�P�m��C�m�M�]
�M��.L�:0���X��)���P袈#n��:�,�C���h�y'�|�ĕm���!�=11�LR�7��)PI;g��m:�?>
ĭ�܃��L��Z���fb���68��)�`^"�o����p��E44��o�3�s�J8�$t�K�"p�������J�4���1M2�;A�ĩ��.��vrH�m��
�������-j����ޗst�5���D��U˺�M5O]y�Kλ6/y�QR��"��S�Q��-����q��+�Yɟ���n���c��`�.�,Y	 ]���s?5�0�T�'&��AMy~Hx��0�Y����w�}�C)��T�q(8օ�`�y����Cm�F5d�..��j���Ď�5&�~Hk�s7.a�399|k+�l����hZJ}������.4'�o��a�?�];��>��Z=1H��a���}�<I�g%��P}1���6x�ح��ƠV �b1���xٻ��h��@�CȘ~u*K��5N�0\�n|d{SM�l�ȱsM����߫;x"PqwS���������_�B<�r-s:
5[�՘1B(1� ���nm�Q�H���ó�Ѵ<���5q�$cci��܀�BsC�q�]����ל��
�k�9@�KM��g^���q<2޾Y��σ��72�cU)���I����6^����|;��ʆ�̓M��MZ <��& ��t�6]@�)�g@q7�{ǸO?����Έ�|�4����C���C�g|�B��6S�\�F�%\�v?��ږUv��zJ7��'hK�E����'���N��c����1�jW��j�����P{0��l���P<}���P�Ko׻�q<ѴGD�.�!2P-J��e�tv������Z8�q�����C(���׷ǚ��%k&�q#�e�x���ۥ���<!'d5Z)@6�=��D�Qn��B��PԜh��A��D���Z����S��q�Z?WtW�)�ݾ��T��M�%�هqW���,C�W:���Et�1]�=:����-F	�i��QP{���C���C�����UC���)n��՘��W�!�7ٹ�� ��yM��>�f1��'�G/3��� ����tU�6s�|��:�B; 5K����P(��{=��G=&� `-3Cʄ 5Bv3�w��4wJ��53��̻��U�<���l����]���`�k��p�
�+�Vc�M��o)n?,���i�Y���ی�� �Fe��4�K�  �+~LG���9:�uaK����2�S]�MfH��Jrk#y���Q��L�3Br�_.�Z�	&T�|v@�� 鬒:�|�(��N��t�����u��|��e��UO׺�1q;?3)�4 AO>����|�F����j*-�����8���3��<aU&}F���Վ�T�f�-�f�皖M�K����F�$���'���\M��>��]�k����KaڟBPۯ�Ae�&:[�ɧ�Ă��g���E�{���5�Һ�_}#�����C+z��b3
/�wwY�*5��B�G�a��*���,9YD7[�!�G��AA�i�_�{�|���4z�%����#=kd����9���XҢY�q��'�|�4������܍�E�����<֢"/V���+�Z��F3,����#W)���yt,�^m��k2(�չ�ΰ��Bb��3��4g�������p���*��ϴ���b[�(������2-���Q�?�c�a�w�~�+'�1� �d���
�����_�\���������ɲ�zv�u�uG��O�J��ʊ��p�HW���&\햸��%�y�1�:˜k��t0�8(,K�}J�{J����-�f�Lq����/����_���xC>85�a�x�"�}�'��+OẅCn�*s�93	(O��?��B1�_��f}���aʖs�8|��C�h-�j� �����	�X}J�N�h+��L��L��y/$,��?�`�!rhO�o;ǧ�꺐ۂ�Zm-1�a��Y�ٌ���w��>q�t8���Z�-K��u*N��������S*��\7Ȏ՘�d�� }��'��*Hҏ��T���$F"�^1(��u���$�x�g-Y�cq�GmW�i%{$���[���ʷ�5i[��]d�����5{�T+������g�U;�B��6{5J��1���f �s�@�}{`��1c��Ђ�o�K��ֶQPͩ��f;�aw�.���b�m����(��'���d�W�G�#�E�_�u]�*�h ��(u@�0Ym��k��ڑA��*p��l����H� ɷs���s
M�~xOh^
��'�B8nhN.]3�6�����r�R��2��k©��M,���*�2��u�����Z��\���Q����#۷bK2�rjqƞ���O"����F�Aw7������p�ӫ�4�G�Z�yL��_����_�&3�.>�ǬZ�ֻt?�Ӭ�R(MԺ騁P�|t���_��gƓ�#�s5��:֘��{5�+�x���ҙ%t��rf�S:����J�z���ǁ�+&x��Isi�r>'����6	�{b���"	���l���윧�12|;_�P+.��>��-&�*�R��J�L���!i�R�|���P�hv�Va�����@D	�@ok:��<b���q駓#�X��vk3��`�R)�O>e����+9�yU2��v�,i�%��r�{�U�-��d�!!�ܖ�Nu!��DD�YoZ"o9#��֦%�����|������ל]4���`�2o�-s!{�9�{���j6��R�A���4��D���  &Kt�yх/���=�qR�yӉ|U'H��x�.�8���[`ӳ����M��<3%�1���+�9�	������b�b��o�����L����*x�H]���)QÃW�~G��o.��Y��jV+8p�&�y�gx���=�˶_C��P�^[��Г�?��"o/�p�j1v�tFe4�B�L
��Y�dU��$3�9�&fYFɎ�A��x۪�����(WUn�t�o�t���GU�m;��m�.�z"�P���A(�
�B5#Z2w��4^Ƿ!��;�M5̹�|�����_���6���+6HӾ�G��*Q瘫�O��*��Pv�.$��)��!*��Z8��~GĠ���g�e�/�w^J�榶���ȗ����F�=YpP?��nS�oZ�WϭcGbΌ��a�
���.4�}�� �p.���{j��>�J�/Xmu��ͣzhaD�dM��ڲ���";���Ә���-Z��Ds%�l�kxpe�|s��d-�lb���K�9�߭���*$�c�l$̷���Y34�0�K�b+Hτ���$vJN����;����Y�d?&�M �¶��w�C�S��Au��1�[1���7���Y��gPz&�M9���/ �Ya�����9y9F��L���Kz`�j��`��L�&�_]���XS1N\��qT�����E>����N�=����s�9ѕW!e3��C�`Y^��EE#��U�R�Z��#}�v�M�|'
!��Q�ӭ� $T�_ ��0q�{U�B��	�9ob�)h�+��1���/H�x[H��x/�E�|�>�zV��f7�#I�T���ٮvDM���F�8S� ���2ى��|]6���r9�7SYI�x��Ȕ�@���N-J7������W
�)�XY��Q��sG�ڣ��T�T�L[".5	������K�vP2wZ1�����ۨ��������h���I��"�2h�>� 1�n|�^c�����c�(�m������@��*i�*�ķ�y��{���*�(���ߪ��M���U|� 6�Or���Q9(��g4}�v%@=�K?=�@@���5g��:L�Qԛ�k����(ȯ�~���D��'�NDp�� �U�;E�Ηh��ϖY���C\ɽ�s�K�.&��,��3T���#�dq�}ݔ��N4�Z��@@���H�oiA�Xa@w��ԡ�c*��j���f}��U�6,̌ ����$�q8p����X��� ��}w:D�y�B����	��Ȱ���l3l]�˖ ��߰�����D5������P���QL�0Th����5�`@�Q�p6��k
%+�Y�K72 Q���&A)������÷��U����`���.��!n�]	p�`�1Qg/��y\�x摝`��`�Ռj[5��p�m-�t�H��t,QL��W�J��T�k��	4x��
�L��������M�lJ��յ�k7ˊX-�i�s�m��;���m�抄8��p�K��a��࿼TP��B��!<Ȝ�r8�o��8>�.d�V����.п�N�
l����^�q��m�7bxt�y���T�K��~L�Ʃ�"�t��E�~�8�n�5.���><%4�iwbxl%�t��w[u�u_�����E��٠�	��o�")|�Sx��^$��8��;ǐ����:��2����n��!�����&�o|�=v;KOmķ��$޵�'f�oY�O=2+#lD�1���lԻv�d�:�&i���bK��G&״�צ����]�=z��e���#q��h�p�����$�]]L lc�O�0��;z�GD��Y����=��T��0�r��5����WX/w�_���;  6T"'�6@^f��3�d�;87Qw�a���ǡu�P���I�t@�Ҩ��갗iw�y�&A4�ҺJc�z〓h�ɤ[���N�i��M���(Ы����e4�^���ҕ^W!�MO�Hc!0�B��XƮB*���;f�e m��* 76�k�����X,�i�yq�
�)B���1��;��R��d�Z�����X�R��jC�"�B2|�3��W$�s��"�BE3��ص��3�B�F�<�T�E���[����ȷ�fj3`*�'ucpō�HK���)tw�4_��X�$����QY��g`D��L���7�PP9J�u�҈c�O�fa�|3�_�M
V��{��	ziS�Y��b@Z- .��25�
�1�c�+(�kvM�1�_sh�W {P`:��e��Ab߅n��ᛓq8�� �yx2�oh�^Xz���q� q�EuĒ?	���Y����&��4`�:��{��>��=��ng��2�"��y�u�J�OќP�.�"��n�m��թ��5@6�8G�j��}���ĐO%k�ڭ�16�A�I�2�b��\�s��<S��J/��M�Ik�6�L�}����u�~�,3d�V�ؚh��)O�,�N���1ܪ�FY6C�,����yW��]0�?��Yv�o_��'թdvj�Qh��ˉ�If	x[FzS�TN)+ś�Ĳ���4� ��K�)�w.+�ұp ��k-��zR9�L��s�b�i��>��������� EM5ƭȗ�IvC0�7�1��>F�!/���O�ؙ{d���׊Q�ka"�=�OO�4 ��>����v��8�몗����u?�[�˔�+��f���\�!'X"o�#Q>c�*̦pN����[_&��&wx��JZ�Qb�TYJ�jD"K� )X8�c_���FC:4q�@�w5�Ml[
�C!�1�M��jM���f2�w�Ɏ��P��� ��2�ڦ����#��׍Z���4u{W> �lƎH���>�:sN��mٵ~�K��UV��q%�A͛��D��L����%��g�4@�-��?D�E?L��҈%���.-$x��|�y��D�����&k�"��I�6U��c��]��<S�I2@�%���'{��4���S O�fӆ�t��Q��۽���z_9m�Ɨs���Ƿ2UX�^.�a�G|��.�+�W!��&K�{��6����m���u��+l���R�c����/�V/C���"�4���>��F�>����Re�<�
�
�^����Y
�a5���#
�q�R���Z���g�$�	m�V��Ю��N-�˶�����%Lx50<�ً|�p0Nɋ�V�^gz�
�����P�����횱�>I,���4�6-�:F5��Mf�����5L	K5��S�K��;O3�(~5i)��8bkf��te�,{R�,�����蹫�y��������@�dw\�]8!t+���KQ͒�ª�<H.;���(;�#��y�	�-��X�^�{�?W��5�H_�a�'aǳ�y�iº���PxY"����}4WW0��d�I>z�l>�Bl-�LO�~����.�ø�,���p6`��U��ԍ���͑n4y� ҄�t)3̵uy�o��x�"F�3�;���o?�����a���D�ޘ�;rJɹn\{G��zj��.��j3x�+�G�����1&��S< ؈��%�����.���i;F��nX/��B��I����P`
�fG�\S��	��o��.����%�Օ�:��������@L6� �Q�7��֩&�����l��c���?P���c�t���
���@4�VQ�F7H���5֧��d]�Đ��^k�(jA퇎�� =��T�����ق��aY��EA
�n~�I���m4�&&�������+�3�<�v�e�W`HU��^D5K��2I��L�4R�R�Z;i������=44P�}?�x�Je�NF-��r����"��u�".�I~ҵ1����I�s�'��7,����q$�{M�nI�G\�wη��p�ؕ�U�/s�M=�۳mq����]	���ː����_�Ų���0�c^���\�k��^���ܧ�����1�.�H� ���s
t�	�B���?rb%���U*%h h��LALi8L�+D6�k||cu��܌��L�tq8��ǿ�I�,�s��JX�T⺛���y�$���8S_<mW;-Ѹ{~�HFE�ڋ)#�'���וR��?,6o���M4��Hdu�o�6�A��taC�Na)�a���Pm%�3�'����N�h��ߍW$��������܊�9���C��J-�`4:E��	m�
�J+��&���ɷKɓ���W��Bj��C鏥���4����'���0��"�z�1f��J�8�u�n���f|�ڗ�hԼ�/���U��㡑T�����JM��ͥ�)�*�J��@�8��>X���E��n.�
	t~ؾv 46��~}�2���Q{�\j�n|O��S$�G��=1�o�7�v��O(��\}@�I;.&�+�&c���/�ܵ��Ms��I!/2n �d�}.uiT�^�a�%�:?���eFOR�?�h�	�y�y1�9�T8PeC5� �+���%�������9���h���Qn�%��L�];����*�FW��\�bd\�n��j�!��Ka3.1�N-fh�3�����j
�
�j����.�_W���*�ݼ5S����o�a;͙x�����$�ֵk��7~)�NNr�E�Cj���U>��V�S��:|8R�?/ �9Q�A�~�Ը֬�ǭ���]W67\���;��C�x����r�J0x��Ȣs3�j��`�9�/�V1�hB�L�}CQ�r�f���4G?�9b b��2�e��A�RL�[�N��_��a��qdC_�	��Q��*ox��֥5�,��""��Zz�pFmwR|�8п��w���}�h����`���m�����3�: ~Qh3�h&�L�!�#�s<����D�ޒ4M&�&n�NM����j�>����}�s~&���!yq{I�?e���'�*�k�K@-�i��$�8u����[�8��u�i^��P��%H�J�U�Fΐ�O����E�eq �j{T��� �Q�{|!��p��9�������Y���3	7˩w�n5� U������*�WldCŏ߰�P�*~�&����v2�� ����B��*I[�����K�4��]#���h}�@C�li��~�����i���W�
 ჾ����LQ`����R��H��We�֕_ڤI!���"�w7?a��<�K��7�)���-��[�u�?�ҽ_2X��(�q�$�Oe�$>;U�p��~��9:���s���-�Ь�y&��t��ݙɗt�D5�.�?��j�6!�ko�=%u�b_�p��!R��<ڳ�!ttU�o�U\�ړ�>6�!��Umap���*@gi�����)]5����p@O<��jlC��Wr2�C6:�g&;֛)�-v�j���tRF4)^�"1`�nL Y0���qL��` r���^�M�~�g��C�lk�����xX�����9��c��V�H�����@(E(�jh�g�N~��D�5��u���_iX�p��=��,�3��1H?�M=
.8��;��$�XJ=vF�Q�(|v���S��II��m�Gb������4����K~r�K�!OIa�9a+����>c��-�xx�n2#iC�}�=�sv�N%�b��{�	3�J�'!?����	��
��1��Qig �jFֹ  ��@d�	��,��:�)���Ê����k[�b�n����D��;,�- ��X"3���Z�X�G�J�"�4�杞@��[��20R�+,Y#n�6�('C�o_:Nϋť�(����W�[�Ŀ`4����ͪ�p@0�~�N���^��܂ ����9�wP5�mx�����t)�KǠ�Py/Pz���A���F��ļ���Ӎ
vO�EN��A��Ta831%PqI1E7'U�����t�f/>YU�X<�q.��)vB3�eqw�@5�h�Մa��:�M���H `�?ҕ��ɚ����*�1T?'s�[���뫫1�-�y�Z!.�͊�D��Cdy���W���>IMM��)+��p�  ��ﱟ)G�i{��^ؤ5G'x�|q�o:�e6F�uZpďk����Gɖ9�[�f�pH�d��k��,��;b�zD�=A+b$�A�+�K+�FY�|�-�2%�坊��PZ+a��H����i{f��'��Zغῥ�A����1���<�n1O�|�0�u@Wy��B,��k9�7.��3 ]�I���p�yx��30Y�IIp
$���+�~�y����n�xv1�x��n�8T�{W3;9D]:�9�Z��--�,�VwǂM����b��z�%wh���],��N	��]�`�5!��_�͈w�7����P�G'kL�yM:�;u���4�s��4�Nr�"�w���
m�� r�� �Ł�������l��#�FrA�-�u�u�(s9CǏ�����嚴�6�:0�W(6R*��>��5忉i;�3�0�����#
�S�\O
�#}��LQ�b�ʑ�
�U@�'��X�	�fS}a*�����u�m��F�\4e�
��� �5�j�=��f�^�/�4ͅ8.�Ui1�#�:���ؒ�dIݠ���6��h[��0��{��*���l��A3#>d����a����u� u��I�Э!�{m�i���8�WԹ@�^�>$fJI&�'�����ēK̼Lh��L	���w����E�ప:���v�h�z���M.������@2�>�5:
����j5���rz�X�v�&���4��j�OW,=b�H�ݘ���b��H�5�@i�J��m���ٔ�?Cg,*un�㔋��8PKI�k^:S��iѨ�k��9����PثwP6�.W�z�Y�{��k�1��K�w�#h���� �0��<c �5	Zd�r��;(^iu�EUճ4��m}�,�0���.(��f�I���Hڄl�H�>��6�*�s:�R���EE�O�ʆ�-^S��>g�o,,O�[������X��[��Jp���}b��؀�N��A���=�&���R%�*���ݰ�$`���S��4p�:_�vuY=<�w5u��v�����2����M��:�Uq��a��G��<X$31�Y	U
�󖕷�=չ$6�4�Zʂ�t�y���c��u&)5���ݔ�S� �Rn��8R6��vK�0T��bVѫb	�E�٥���ٿ��{GA����0�ް�}4S��6�����ԣd�zL��2͗��g)9�qT<����ʋg%�-S��}���!/>zҤ���a�o<���^�PLw)t�t�t?����K��7�Ҫ���(�?���wv1U��o'�����!x�������F�$!C��ۻ��K�0���A5�΃��3zO����W�W�,_�햾��FȦ7F)����\�?�Z""W,?.���������؁�MፆBx���Y�Ó�˭�><��C_&R)�| Ɋ8��Έ��NS�OY�� �I�!��y��뉝ۅlA�9|�&��#݅��E	K��ic�*��Db��9�.�oX���t ������������xʖ����|�Z���m�Y�m}��/�%ӏ���w��&��9gB��U���3<\-aS�u�1չ~(�J��X��C�˰�o�i��.s���E�|�[�L�%�w	��0���ߊ��w�"z㚼5����:���7���E�'D\�z6*�B&-y~L㴈�>�?��G%YV����2\�����:�I���n��r���+r�;�h����c�v9*�h�>5���|�[��d| �f;vR^�)F�}��`���:�b��c6G���[�R�d8Z��SD�B �2��,K�D�s�@��Q�%jA4�q\��ݵ��X�/��D��X�i����dC1��H��a��Mڦ*(��Ooc�_�%(lpX�$�>�rVE�MQUbC��G\HV��)6������PV�G���}�4%�"$^J�/I���e���^e˰�V}���&;*��{1�VQ��jOԟHI�N<��h�k�����yH�T����������"��*���H*x<6ǝ֪�T��������"����)C��D�p����&�3$�S�aZ�� o�J�X����#�c.��݄�j��L���/_�Eg��j�q1�I��W;5�M>��ƚ�*o�''�ॿmd��e�;R��K�s���5��I�Cq./GkW��f-2���a��i87\�p�@���?�����RdOs����<�ya	��<lo@�q�0���1P��Q��cQ�l��d$�t �vD��XzP04D�<�'W�gO��(����V/5�(gf�I��1@L��֒��%�,'�튦�PS~�ލ�8�Ch4z�$�wC<)2W�G%��1)&��舶�&i;_rG�{>��H`<���U{Z����i���SN~4����?�"3aM-le�C�c���X1�`�m����d�𗋲�Ȍ؈D@�-_
"`�ۭA7������xɶ;Ҧ�'e1x����Y���Dr�-г��:E11Ҫ��*�-)��ĕB�$�lt���4�p��1�_Z"�� ���	������ �7��7�Pv&��@*g��6��1)�$y�X��v�߅��FsU[nw'�a���Bކ��p���_B�e�0<� �x%k ǅ8�m��G�M 8oem�)���P��cN`��`z!�{�$l~ߪ�+WE/.?�7QF��	�EK}�a��-24��[(��wv�Ao���ۅ�Kb������GMa�+�<���|^��q3E��׸�  z�W+�~�q���'@^\6u���О[�?�Tf|$h:l�<۶R*���^V�r�rO&��1 � 9{*�=�YZ�^�[�[�e�	Ѓ��	#@��F5�1%UT=�p�TZ#v39��a�5�1m�KJ���1m�r̎���s=��Gsg)}��'�z�_�v�e�QGuK�C3N��O���7�ͤL<e�<o�gP����@��<T$}���?�8�����-!�(?���#���GV*GP1�*���s���rme�CXcV�b�/�E!�;�`�M�)je`�_u7x�QU��f�E�k�k���D.�3�PH���;�_A2B��\��ͮ��{���>����D\si�<�5�����N����r=j���,D�!���}��jg�����T�v��[� y�ˁ��@APw<�>�?1���`g"��ҋom����
�cϟK�MZQ�*��.z�5p�$������6؉W���f}��+��}�r���G�h ����N�z�C�q��Q Y�U����a�O�f�^q����k��yA������I���
� �,9 Q[ό�:SƔ����C~HN�g>�x��]2��S�R�`�1��LVF����!bА�2%t����A]�ˠ��4�@�ߘ�����3��w�"J��W�5�,��
��/��P�\�o1_k�h�_N���9kq��}�j>8s��ݪ�*���9��e��v��Q���Q�1�s�˹SB*���ԫ4�^0�7��M�ū�\��{����+s{bb� L�{
<W3���<��C}�g�Z�(yyb`r����K����SfN���R����)���9"��]�%���@G� F>��g`���) �B�h:U��?GӜ<b�'��Ǐ��"�)���ۂr�����D<��i@�s��|�q5��3�BnFb=�O����r]�kZz)�y��-!�tb�p�V��O��`O�����c���+>��Q ����lpc��[��r�7ㆹ����H	)k�.�p��#mr�Y
8�W)cUbI�-Q���)�{^tWϸ�
�E6Ѣ�MQt���?��t��u ����Ї&X�:K .~DA/P���Cx��}�f!�{t�{��%A!@�� �%��jν&.e?h	Z�R��i��:��*lO5@K���Q@��Y֒�_Z�.y����&E�π'��s�(F(�6q��W!��?�Bz��?��W��@S�	vW(�����?�K.�(XM�e�d�xvR����l����p.S�8d�����s��Ad� �.֚�NOd�_9$�b�����"��6�DE~���1S���c�p[f��!���8��������Xi�M��0�O�dv@v%�+e�J�L}x��A��+��F(�e{"���+����E�Q�����)�\��^!T������*��g��8x��;Uf���.�d�{m���b|�Vl�3x�u�eԶ��΂e��WV����CX�֯��}��0<*غ�����v��;�}d���)���n�a�-���O_ ��������ߞD�tF ���h��'�7�"���	�nu[R˛� PO8*�=Dv�D-]|p�����F�M�)�q���g-�������"����%�{��Ţ��y�H�nɦ��m���B�V��uΏ|�\�S��U�K��x�Z5dM��*��*������E�2��K��+��%�t���(��g�^!�V�Or��� �o2y��I�킱�����`Xi�CК�/k���f]�P��B�b��4�$1$�m?�I����A�a�B	�[��^_�����\7�B9���d���)?oZFY�ػ"%|Q[���>ef��x��b�te��t�ߵ��9I�X(�����V�ls|&�I�-�TX�֫B���h.�`�4q�U���B	dNrV_sK�Ϣ�%�9w%	��e2�&E���k׍p3D�Yy�>�P��2�A�CW����^*��`Ô�@�
�\�S�x%'��N>���~�mo��rn�0��m�xr
V�ִ蜚>A�m�s��FG'��-�{%��5���"���r�����Tpe��rR�E��?�}���T0�*��^�z�h�����0����
-�Sq�k^UT��"�2����_�Ktu.�N�c�*� ��4�w��`���K��?������Xנѝ�	nUt�N�ʐ�1�����7 R�HN/h8Q���pRK�]���+���X_��lH��Xϣ��;��M��D���\�,�"���"Sh�$t�\U �{�c�̋mՏ^ˇ��������E�\4z>�(9�њ��Y��tk�>����rȈs��>�ZM�y���3��I�|�$J~���Vh����<RUZ�����T����9�%�En�}�1�W���V������;���u1�4z�9"��3�+v�3m�!E	�1�$>1ǰ�0_9�kԛN���2��@F�k��k�k]���+�o����L���-�N>��,Ǡ6	��.ו�k��x�[��P��W]TG���P�v����8r`�����.圛�ͬUO�G�厉AϺs��,C�/3b�s��y�o3C4�XR�n}�i=ɛԪ��K���o0Iw�ؒ�����0m[��3~o3�{;�ad�7r���U9|^�Ҕw�����ɥSC�8];���h�x4����F�V�(����\�};N6	߇ŉ>��B+)��r![�J������z^��H'�,�$?*)��q_b���-��`U�(�)��m�f�s,�3����d��f�r�Ԏ�J*UG����Fi���K��H�K`&��� ԑ,�����v-Vj�7�GB�^_�����P��c�;0��P�aj�sЩא�������`���_��j+Ǖ`�B���#V�,}�Z�g�j/�1��2��͸&24
����R������#�]�Ԏ?sϴçnPd�*�i��qv����4��6��GMr��8���|�~W���f����3{(� ��-����kD�^��a����I�L��!��Q=�H�Pkg��F	���YINgA֞�4�gm��{�,����S�xi�_݁�l ��{%B���͉�{���es{�ڡvQ�E��p�r$*�gQ]�9x @X����c"C��J��x\��p�R��z�j�:���wrqh�Єo����u]���m���n�!����s%�V u��55-�l���Y�89��߻�a���B2j*��"�X�1�1��e	̧������ ��Cq�y�.T�D^ �6R����Y�Ex��bY�3D{�o<0P���@��`���j�|�yM�7��F<�I=���ǕA �~Z�n���O��{c�A����A�x��3�\�G�@�k���'�8Y�Ѡ	w&��\�[8:���B�Lz>���F�7��,*OYѰma3f��b���?�"fz�Hy5m.�c���+�N3���^$=����������{U'e��`��eI��9#�-8�&�)y�ܹ݁דEo C}D ����ό��(j��c��y`���͹��8�N����<�L� 8'�d�>���&�8�b�HI	�o�C�X��ҁ�+�,���!a�"7d��]yE@��]ۘ�&�M��AJɲCi�c����;�n�cŷ�4�/H�^q����70������88�M�.��,�[��#��Pn�m��F�tpY�d*�����^{8(*���в��˦e-^	��\�P,<F��Y�y��a��) �;�>�
�鹎r8<o��C#���ÂRC��X@O:��i]���T��^��@������8a��0#b��ƴ�F��� � �M�P��������.O��:v\��O`�����mԼ� ��#ᬟշ��@��ݏ��;Z��Q����KۖO^B/�E����n
��o��<{�C�O���(��-��ܽR@���B�FW�N��z=����O����K��ǖ׬__j�Ӂ]���AC�u�*p�Y	�B��:OF�,쨱2ǡn����TXLDn0�c�*3YG��� �Ž�TSq�G55y�q��^�`��^��*�*�?��w�m�֑l���tj\�b[�1M� δ힨@�A�&�Uro:zh1Rg혠�pk����X�\���ҡ��c��H-&$��l��%�nv�R����u�K����dm#�M߰�j�Q�&R9�V]S�I׷��۴׼A`���/ӏO�8�2�F�?T9ڌh��c�����*���";���;x1����q2ч�I�|���!H�������<����U����!�Z��N��\D7���MM�(g8�F�,�)¼��+J���& ++��:���|�a�k� i�,�37�����q��M��ʘ�	l��>�c��^��(�b��ȳd�����t.�=6�A٬Uղ1>��rK{4�դ��x|!m��R�<9����# ��k�4��rF,��W]\�V)}H��M[Ț^3�f:?$}Z�/������-v"�����=~�d#z6�xLO��k�O��F��#g��I�WU��`7C!��~��k�B��,u!��:�BΌ�.���K$��N;{�8v����Pv������A�ihʧ�'qB���&"kJ�XA��u�GPz0�ծ�է�1@M�r�N�-����a�t�t"�&]����׏wO�W����������vv��u�vs�����-d��fT�]�::��j48uZ�I��|EWb����v&q�z�yK׆v����=���"DmR&!�[�q���=�/@Ht���!V-y�`�q*)S���Wk�Rv�+���������m�Gl�s��<i���5�GtT!3��Z��C�y�۶`�sF��h޺�E)�$yo�d�t(F�8}eiB�Nv_�Y��ioZd�(u��_��G��r���
L���kyO�ӽhX2��^���y�Z�*�v�i~C��.�<����l���:���z��Bl�u�2�~�{�Vp����?,8�_GE����Q���4f*��U�����=��px:n&���� ���#L������i�3U�f:�g�����}I���֥�S��#'E"R��eh}���՞��] brР��-�r��d�X���e�8n�5�U_>)��_�$7�y��vB��N�s��_���Rּ�]���UP�����Uv��D�_Q�ZO08���e7�W�.�nmv$t秆kͲ7�Gf��>*"�2Y'K�x�qXi���Վ9R0hq<�"�jLh��ʢMH#�oiz�,�Z�c[�[���nN)�#��9��dj�����V�}�UB�/63fYB���|n�c�]�;�����ҝ{j�7��3fVSnm.����,���A
��>����OG��=�e�AAp?�����t>��h�p�1�&��+�96x�&|f���7����J�B6ݡ1Я�����V_L�5Tq�[N�]�^�8���t��*V�����y$ȯ�*�k��i���#�%�X��+��3��K0)�Ͳ�`~�zsB��a��vEQL9"kP�(D��"7vr^��qa�|V�b����}�#�ɒ0�
O�JJ{=[&������5�����_S:D�NTúI�j�H-CeJ]�id�(N�Pp�P\��#�{��S�"�4� YG|��ǒ�̚h�}�8�c��_(��1�z*|��p�� "�«pQePi�}\�^:�,n� }sr�^���K��ܖ�^YCwV�'��A;�c�&ǽ2*=Bk�J��V��ն�����<`~�S�ɓk&s�xU_P��lW�l��/C�;}iJ2e-M�)X�X/4R����|)Ʉ�{�w	�H�w��nd����4)��y��h}����'��
1��%�J�!�w�<:�}��*���e�7|nM�b�y����;�{�����`3�߻X��#{n ACy���\ŃL��$a�C3�KA�,�
`P�u���E�W]��%p.��Z���.q��.`���y������[n!��G��Jj�����h��u^�T��t}#	�a����d:��+�.il�9/�k� Ѥ*�Vz��ګ�'WY�:x�8������_�#��mD4un�8���O�ao�3��_x�ڌ�l�[u+�v���v� v7�Hr���)OG4��R�K�1��*�D��~J���Y�h�����|Y&���~r��q����3 YG�Y��y�_�	�)��u�J�6*���
,�Ґ:+sT/g����@��ȝ�q�����`"o丫 ��8�Z́xu0H�`�)W��Ahl�&�Rt���؜���P@)DNo}r�n}:Z����q�7��U��9Q����Q˸*���=ֳݮ�ϕ�E���f��Ș-�ǅ�*G�Ed�to@��@�r03�����9� K�2nbKTq�"6ԥ�>�|�J���C��)��8�|J���Cm����!�|���Ϯy�s�؅�Ƕ�\���Zc��ChO6��8&�k�`��29Yzb��7<?N�(�i����u��+7��d�!�12ex�����6RX-�0����q7\N�B��ϕ�C�7�C�uX!I5W-.k�g�6y�%VQᨙp��q��R`h��:�ܠ�ai��?���V~9'���7�}�Y�j=���
8Ep��q5AhIj]WFC��������<��1�H�K?��x���e�p蜆
�l��`���(���?
����B�.�}7���D��SP^<u�7+�<�|�\��8���������:����V��3������3R��t�j<Ki�x��^�6@�hW�|��y��=�rq�uwkO��������W��ѧCXtmF��{��n�K>^�E�T|��������?;��)�i�H�n��[l���&d|r�����b�T'��[յ��vk���c���Go�`��`�6�1�wF~���zy�&D	��NɁ�t]<;������E����SW%Yh�����U��0㮞�+:��㾌,#�� �ׯ��t�}�}�w�Kh�M?�E��g�-�m������5�	�u�j�'og�>m�/G۵��uν����;~K\<8��OMb�86(d8��3�����$~�}Q
خO�/j�����E\({ȲV�>1%���d1�RCq��	
��N��H���2�N�i� b�]����n���ۮefQ/�Ss|�C�@ы���	�u���R��0RE,f�o�"�[�2�i����J�ۭ$3��6w��L��<Q�kR�X
��c#�M��rc�ˊd����]�iPף�O_��W;�y���Ɇf��L�
�����>�����
1$�)y�&>IED,�Der.�P��kf�鉶�b�d\��/�/G���j��9��q���@��������"Q�f\��6׌~����p����.5BIT���0�Jĭ��(� C���n�&�S,��䴞||[[�G�������4��0��3�$��M��+A�D�g��.��<����i�5�3�Y}_�P���ݯ�3���N��q�nm8F�
 �PsN^�m���4��R��"J��?���t�0��3-=��B�����6`��-D�]��o�)v�k�I��@�A�����h�sF�Y^��w���-� i����i�2�b�b|�fȩ3�+�~��	l�<ήX��
�f�,�'g���EZ���uZ��@�:~��Y�s�O�4&���������i,��,;ʸ�j�4!�I�/��8C��f_�%�A��$�t��K���&h�`J���rb���E&���[��Q��:t�m;�嶫J�_���o^/+�C)�A��b���[���Mrt��b�̘H���Rl$�̬�[X�}U��r���4[�9��kK�j��������"�
ն���>t�)�L�2�S댖�a�,sg�N׮0����G�w��6`{L�5,W[���-��.���qM�>�)D�3��9}T�(4�sL~&ȟ��G��D�7���C��WG�~ɁQ�!-g��T�r$�M`i&	�Ҕ��8����\��֐be�Z4A<Zk �T����`TĀj��������^9֋����{��Z]�2(�:AT�Sߝ{<�r�h2f���(�d7q�V5��؛I�a������.��I������yYͺ0r2E�&8��N��|~��\�9e�5ۘ�K�:���ʢdI�e�{��S�����&5�(Iت����s�Ԅб��@}^"���Lv�<5�����Ƿ���U`�0K�C1�8[�{ $��5k�D�O�a����x�_�'�

v.��9̬D�g���O9�C�y\��
�Z�. '�ޞl�-���\�*�Y�DE/�Q�7o�9:3�t'K��Ȭb7���O��X�Iy<�kf6������ƥ�Y��=����K)�߿yan:� ��/����th��|@��I��o?��\s�;���������I!;���սٟ/��7�f7��y�s�o`,��	}B��~��!��',-l���A��W�7�ḑ���=l֗j�t>��esF����J�0}s�p�(X\�sq�"�_
N��ꐼu���V��5���>�#� 7�X�V��L����0�"(D�>r�4@�V{�Ah�>��k�`��TӃ����f���:�d����8�N	O�p����|��\����R* ;�tZ>Z۹��R(X �//�ێ�'���鶂6�#$pM��0��O#�W�mstc�M���Y.�ႂ��불�4���Z��K�c4����T�$M��I"���a�Átx��+\SB77���������|���;.�|�c*���P:H��xCrv=ѰF��1{�K&-	u��`rX�����`J�U�����-�|�[<��J�XÇ�M�g���H�,����@�U1���Hr�d}Y�*0�e���A*2	޴�OQ��w�Wh"�����߳Ħ����ʍT_T��ͨ7�����56�N*	�1~��S��r�,i.�j]��LH���lH�4�U�h)��&��g��[����;��Z��Ո�u���B*s�f* (�u�0�o���O5LL omף�=b�Or��yN����gW"�Wy��fY���Q�����m�u��O�hc�De��ie\��4�t��`�Ď��|r3E5���^�Z�M������%H)�vB<�����a�h�����$�nX�L�>�NCh
9;����\h]-dv��c��'w�-��-�oڹi��(	ez�d]Ĕ�s4�~��2(k;wF�|u�_LAg��O-b�65Ԃ�.΀g��Pd ����λ�,�����[&����].�cȻ83��WNG��j�n�QD��+�ī��kոi��g�5C��z3V��O�V(1M�'��v�^� ��-��R���H)�h�yl�@��DoB����hb�M�10-y��i݃PM7��Is�\�$fd��rd�	{�'��0 6�_��� �n:� V������ �{ 0��W9\��>w(R�e�'�Ϡ���w���7g� �5v����ſpLY	*��Yi!�<�2��|��2�2�AA����xl6p�5��W��Q��bR�����ƿ�Om>z1|;QV���}}~������m��+)6��t�p �:=�ء�=J�
��:����R"e����,�}_Ɓ�N"����'��\��|FUq��.x�L@��̥���7�(/��{����4}X�]��t~<��G�SS4.N�hE��W�r�A��ex5�E8)29*' ��9Jb�%�*`�J�����֫��:��PgY˹I·�M�>�>r�rW�z%�V�8�������ؘ:Y��S"d	*�~WŨA���y9#����JԺ.ElΩ�^��kd�7��RI/�j\�Щ;\���hj�?Q!��T�h`��M��e�{r����=�n�X�p2W x���!��0��i��Z��i��" uq H����O��mv���d��ӻZz�k��X�=.*�ֱz�Oy�%���*㉚&��l+k��!�)�7���ؙus�J��|Zd�dK ��ka#%-�܍o���tt8�0��T-���/I#3����c�ճ
֘C5"9j�uWt\��"-_N�!��]1c��L=��&�m�^�4��0�.z���gG4Ko|w��������a�45- 0�j1ϛ<�	)-~ ����9�!��< $���D�I�����a��X���|���Z��ō�&u�б?f��Ј�͜e�v��7=�2U]ߗP��LSE��H��H�8����Z=7����>KS;����uݫ�c�%MXY:#�y��|���KwO*�Ȯ���.�,�jB�v[1|��Tw��������wKX�!I~��@.q�P�B~�����Sڀ���=�3�K73�d%iV*4�h.RN�d�v����0��wHYN�r3Uy�����߂"��\aF}�H��pAk�F1g{PPaW�Nh\�����<԰Jg����vBe�6�aV���S:e2�[�K��H�/0���(0�8Q6 loO�뒩[,e�͒�e� t�D<�Aq��w�~�+�<��)&[��3ܟڑ��ЂL�
#Ѫ�;;��p�B��Ÿ�հ�DqWM>N��M��t��F���ڀ����焭�|U��=\�m�Z��.c�Pr� p5�-}�`�6Lk�g9#�M6�??�S�d��qL���^�~�ƥY��v��o�pӽU�%LOHL��/K���Q!bP�#��D����f9&��s��|	�S�{�H��4*�>��[J;���Ԗ�&G�3n�WXp�zy^+w�T�b�稚�^N�N�ʋ8TN�9�����.1�#����t�MH�l4R��C�'	+7V�m:J.X�N��a���o�b�NL˝��`��\�H||ꦏ��U��KŜ ���Z-�A�8G�u>"h��8Fej	���@/,��:h�wF&�E��y1s��I� ,L��*L4��Q�ئ������v)J���A(!y(��3�#q��?ľ���(�Ϛc�8�
%�h� H��#��jO(R�<ǡ�@�Xٱz�[v(�<�ؿ<����1�%���'���C�6k��RQ�C��$�$��}nN-��B.g�$�����Ԑch�����c��|��!Wq{C�D�ܦk��� �>�C�}^b����ە�_0G�7>")Q[����T��F�h��Aʝ��� ���f�s>�{I
I�z���즪���CN���nz�۴��ռ#m/��l�4N���(��n���EQ5~�*�2��޼��@��T�&^�*l�G�i��H ���v4�W��>��pK a+;N���j׼3�ӛq�Z4(���Д�U��EM[����>oï+x����Ѳ1��>��{�5���ɼ]��������~��`{��༷3��澫Lc�<R}讵��7ö��y~L*M� 9�,�A�e�p6��TgY���݇,(�gbm�8�� N�"�+��G�L?E��_R�N(I��U�D�+��d���7��-c���Ϡ�z��,hj�0YG�;��c����<ז�Jұ��o(����]Ì"і��ʁ�'&���Ou�۴��Ț�6�o�2 �'(�E�{r�g�J�� ��܆�wJ��q����GB�{��{͙��<�Ʈ�:2*j���ߝ�����~پ3�F��� ��T4�Sč��I�������p��2��J����P���,���4��U�k��L���+v�kK��e�E�R�e��H�N\ ���@4��w��� J���ĳ���iI�??����+8�T�" �}&\��Ұ�4D��5F9ޟK	����4��i���w�̳wW��>��X������Z��x��=P�� &�*��Ƞ�lU�(�N�x�X�օ��s���j~�^Q�@��:~�؈A��MK�գ1���m�� ���z�8���_ĝ|5-߫���ŸN�c���I؏@�$L�5�9�WA8O<�M�D��!`9�a�o����o�`�K�����G�lL8L��R�;�L#��H�Y���ㄲcX�@��dh|6K�%���p����r���+���O�g �jQ4�όq��;gY�-�o{ð?�>}1�`��㏈`o�C8��Y(.��,�>���qi��ʚ�;���	=	9&�Hdi�8���.5�ci!�� <n�W�[�ɖ��wG��3�ڼ+�{si�A�0Zt���l?�����%�Q�T���'�6|@��HF��˵�I8%�< <�L��C'?ܿ�C�0�(+���;��B#��k�*
}��@$~bSߓ�����&�]#�˙,��*&L���q�PA��Yu���>�^c�๳���s|�:�Y�"V�^���db<a�i����?�x)<\[�_�=�/��~�pZ���<X'�x�Aꅒ[dƐΤT�ޤ	��Gŏe�A�S[g�q*�p�MU�\�y\<Pp��'�SX������/+���hn�+�d��`��4X5yI��/��
��k#�V�������S�1Ѿ�l���;ަ�O$��A��_��0��m)�(]w�������ջ����]�t�~:Pf@�"�_�Ә��'��NH4Ԑ=ǲ��J"qJw.�L/�\5�CP�H�wnF�"�Ot��*�[�o۔;�wzۜf��k�����������KZMh�rb����M�uP����}���D�\��e`�Ǝ{���a�x9d\�W�����)�$NФ��ۑ�Z�5�8��H����dTƣy��VD���G���� �i<q:��!��n��£)"/�*uRw��n�h:j��w�սVW��+�L����7d,�\8��\�r]�AQ۩Z�١�g�w�K�P>h��x��O�ǣKʱ�<}Y��=˔(i_r|���N�@R�S�<?�J�5�w�ĭ�Im����n�%0/:$�w.M�4V�Q�I�'?M��{fMuQ�d��1�6o���@ea�[��uD���.�}�&���)�C��X�1�n�^�3+!�ևw�����m�16p�̀�)b>HG�\{�9Op7a�4���WՖ�vD�blCE*"��P��g+|qʜSE�Y�+���!���,`��(\q{G�GH)�'�K�zz�3| T�KE��U�)f���D����%rb�և���	1�(�;�J��",�yޥ:�9������L.�-����B��:��,q�G:JY������ĥ��`�Wlߪ��d�Y2X��<���[r�����Q��܂Vu�y��@������Y�_�[Ts�;x�+�c�a����1�
%M��疪ă��t#d�q=�=F��e.��_$S_M��dq���};���C]d�y�W����HT[���4证m;��	�����i�؈N`O�5I�����.Uh�*��7���S���[�a�.�Z�΢h%�7+8�K6S�����g��zȎPy3d
�.� �4[Y_3�����
4�O1R�j����s�
�{�׸���U7Y�#�H��8d��H��ʋ�l��E�5AS��~n�{w����
�$��4'�o��uq��u�&�Զu`x��0; �#�T��y5�����U��zZ�����j��ׁ#����C��i�~�����s]̀�j �VeR��e
�����L@�<t�p"X>*��r�-&��Rb�Z
v�ˢde�Ohߔ����ugE�G.q�Ϣ��3��=P��~比VR�9ڻ�l���_h�vq�³��d���1pr�'R,Qh����@�Y���#��M&���*�:b�OIU�5|�/ .��#�PII6i]��Nͧ�(�;��E(æ�ϰ�P_8%�.�n�o�P�"��CPyq:�b�Y��K����J,��|M�&���p$�gS�t�M�	ں�,P�I�W�$����=�ݬ��1���]��$����OИ��"����&ig4%B@�HB� o�����V��9?��v�
4H�8���HdSi�?�a���X���Ɯ�y~>��^�|�  �o�N��cF\���4U�n	�И��g ��|5�ޤ��?�3k%�[�y�{Zjϧ��[VZLF���'toQȨ9�$����zz�<��?M����v��ֱ�4fq+f�_b�Y%��� �L�h<�Y�mz�&y7��M���~�� ��������x͐�D��
6{�aTH?�g�p�<���\t�)P��@�۰�J�������B��Cv-GL@�q9�et������?k������bgX_���<ʮ��S Xm�$�q��-��ܑ}������JGk�ئҼ7��e�"�D�.�GH�Z�r!��qi�f�<�N����T�����3���7)fHG�~��2�]�A��dPN����U%J�Õ�=�m*.>�m2�@��ԯ�8��G�������s�p�
�
��#94e�o���d.��i>1�����������&h?L@)�<`e�����}��딪�z�v��ɇ�GQ�d�^I(�q��k��;�061*��.��'Ȍ�� �q%�\�NVq����(l{��9�e���(F��km�%������\��f�+̵�UifR5-�;���F���bK������Q�:�G�8�֢2��ˌ��@C}�Y]d�4V��0�Z���.VȈ�b�^ ���^�qk@˷yv��zm)��� u�$z��>ۗ�=[Vz��2�	-������Td*Ғ�R,L^E21Q	�5�����~��)'�q4%�z���)u���6�C��]�RT^1���6��&������<N���
]Qk�z�8p>#�4���S���Ao)9?1!l�(eU��uȾ�K�y��pD��(Xa+���\�9�#����O3"�}q��u1*(	�J�o�*�}lV��a�i�Ag{�+o_
�j1��u��*���7��8:������N�)ͷ~�g�m�K��]]�H��1I{[��SR��W�	�3."�f � �e�u�J�`	���La�a�-I�1 ��xk� G�ٿ�]�Av=`W�q-1ӡ��G�#�^ ?u�
7\p{|�|�z4��vnǩi+\�Q딪���j�z4�8QZ����"�9�-�����/�+�{cO{yc��'y�b_#A-�OРRі��F�dY�T��K���+��lwU��a�L�=?�u	�۪�O� �<���	S1��,N��tSHu���ϐ�trʩ����3�m�Pl�s$r�L���Ԍ��s��	�T2�ӿ��*�N����M�F�ays������y˛-�H/�S�4�{E*V�U���N��<_$���-@`�C��ΰ~��r��%9���n�T�j��w6���/^��;Ĺ#@�gi�)+��`���?o�Pq�.ci�ඊQ4?�x��M�3u5�ʈ�_]�tZHؗ���S����d�O� R��<b�}j�Ó�s*��]u}��)e�]����*`l.��
��*՗|��B͔�ȮHA��eCn�E�7z����+���:���H�4z~�M��~�)
b�6|���a���B_�4[�:}�_@�t��rf@���9_V'�����}el���oOUݨ2����nʑ������V�����׃�q�A73�t���`��ėRn�3$���;z�D �լȤu�����Αf�'z��<%����6�i���Y�t�*�1<�m_��Gck���� k�;I&�YsJt�7����{���3�&D�;
U�ڬ���~��1����砩5�j��G5:�s�"�>ࠞ�G�7F��4�Fv����A�Ty�JWC�eq�կ����C��*�@���:�Ro��]UVL���(͈x��χ��ʴ��?�6�%g��}+e�r��YR.�ha���ǋ,�>2]��"M�e\/I��>��±�+b҉�G�	��3-�S�=S+԰�(���
7 xV��oޣ�<V��H�:> q�uO���Z-�˔"�k@]M�R�H��y�ئ�PYKȈT�-5eK�ɏ��ɲ���7y3!K��>c��Hb!�; ���Z�p̕��1y��9�R�%�%�k�F���.��פ�|� �.�0��O=+����R�����5�>�8��K��2�?�:ip7o:�N �'/y��W��&iη�:�����`����R�Z�l�F�g��f��p��74̎��܇a��0��\o�>e{�=|��W��p���|d�>�i.ؐu{M�EF��n�-�}nĩ÷ot���P��[�n�#�*��2��Pa�f�ú�nYŋ����tse��Ǉ!q��y#�G���*2�8<�yo63�c_c3�d�@mc��bL���ST�C�3�k����z���J��i�<��u�Ea>Q�,#�G죭?�ߘ�l��	�I
�H�f��@^���b�{��:_��o��� ���K#�^�Ɛ��2���S�6$�aqa�)ۛ��}������}��8�xT�*]+bj[ń��{z��{:uᆀ���=,��x1��Z��N�K����ިYr=�0�R�G�h���HI�r�y,p��[~��"<� �do��CYY4�g<���n�Jiܚ�vs��X:Ѭ&�x�vI�D
�R0;[s�|��J�	�����-�	��R��Q��`�"�+r����;����{� Р`��2���o���,�#G�'/�u��}c�#���J���V���4��Z���L���\�D/�@�a�Ⱦ)�?�%I�N��M�Y$C[��x����Y���ſi��>�k��$�G����%ڶ�6���/3+�p��B mS�^�-���.q-�_-1��=Sw`�b�J+p�Z]>�3��K���ftD�<�(�'����4�6�a��~�y]`t<�Wz@���8��KG� �LN4���H���sa���2��d/�?p��j���7y�,J&'ITR����_��$��V�������۾Q�L��95Z-���@4Bc��Q/OP�(�#w��R{�C�h��ʵZع ��b�_ax�1�t'�c��6O���+��;��[��].���M��FYB>ԈMy_>������M̂(����1��'���5!�w������l�b�ǒ��"���L�����Y-��]�"��\�G��3��&䞒OV����.�G2ԉ%�%��;p��B*⢦��r�kS�LV`�"�/���� ��l,Kk=ĵ�d��ִ�f�]	�Ka� �-��~���`-�9��=�N\��֥;�9�/�_z>
]
� �f����mB}qj,L,�볰PN�Qt�t���;�{([ �1w]P͟��JHꀑ�V�aD%BQ{�c	���NcƗi��S%Y���GvQ	h�����[+��L�/���<���u�������!�8]���^&�M2��h�[�p��:ǖ~��!hT���~0�W�c!5�N�'x�og+�i���H@͘3=N�!L\��4Y�O�(JC#l�.�шi*��hy�ړ��a�!C]'�z)����1�s��1��qv�A#�o�h�u��_��g�C!�4$��(8�n��Z��ز���B�A�����U������K���%O��f�!���j�eq����)ڷ���;�g�/#���`A��U��Vq�nmX�0�)�������XWU�O�Ck-�߃#�^
		�D?=e�Ǐ6�q^��K�*�!���Z�r~x�%܏$��\�[�17��隥>��23��uV�Oi~y ғ��Be	sʣ5s�����ͻՆk�S��G&�]�d'���$�p�!���2���K�K�VCu���#5���͈����Ą��h�����.:�lVu�@"u�w��-�4�_���D��@�Q	�;:>�}�}��_��]~~�镬_�榅��>~F�k�{��:8��~�mM����F�DX�N��xb���Ђ4O���dA	�	����?Tm�&�ҟ��w�G6A�/���u�;�����&֜��*�������>��Ǽb�g���a��(���戅��J4�Wz���_����4��L����?m#�Ӵ#u�ȯBP��X��B���2cݕ�.帮�۷ɖ�8]{ �]��U�|&#�.^�E�'�:�7J�2Y�y��ł�'k|��w��d���B��S�G�L�d�{�y.	�s1�r�I)[�刊�|e�Dzb���$���IL#��[��`�<�O��%���]=p�)��&*p<�;���  ��x��غ$i�p�Y����{��
Z	o�es���q2o�ۄK�f2���>���/i�7�4#�m�q�/�jɃ\�r��@2Po p��],[�@���R5�e�dř�BI�pt<n:J�I �����%d�!��[�n�d,�x�2`���Q)����#f̔�o������[<���ڎ���h�$x��ً�X� _���wJ�v���p��C�CRa���a�����?�R7:�;���o_��,&��n[���0\�h���<�b�ךg-F
<)�Es��\�P:]�_�shXӎ�,�Á����I��5�)e{���� ��5>r��ku
���U�3��NNz6��9������>4*�+�o 4g��9����$�$�z"YCz-�Q�xS� ��Vұx�+@W}�i��1C��90޽�lq�1@G� 0���BD[}a@!�(o]����>7��&��!���$�-(�f����A� @�K�"��#���<�d]t�Y��v<一T~	��EZLgϿ��f�/�>k��6����#/ι����aU����g�N����B�wB��K�xQ&�,��&�=,��KH
=ӕ�W�O|�P�=���8�[-�!q�s�֔�?�}-0�,h�������N[��"�#���K��mY��*7P�A�ݏ�U�L�L�ٷ�X���>ʟk1B��EÍ$w�\N���z���qDw�����=�1X'��¥uE����	������;���3n�~�rЃ�+6ݿ���UE6,��C����E����5��|�s
�C�eJS�Ίj����{���J�"u�ۘ]�@��V�}$v4V��ք�lC~�)bi���dӾ��[�3}y�C����Z;l�NSzC㚞":�ްL����J�+�zZ'�pz����ry7{�Jh0�~���"&�d.:� �tP ̇��ӻ{}�������Q�o,�^L؟A��[a=v�Uo�t���Uזh����Y�蟰T�6v���8���,> ��2�� ����>��%��r��v�sJ�k�(���I���O�s�_w��r�a�6hp�����*N�Є�!U�D(�J �?�\p+Y�Q�E�qM'>�]m��
����Q,�$1��w4N"P��c�v�}mW�-$ބ�ytt��l1���f�Q:�
�f2��E�� ��b��6h���+���"�T��҆b����l��']�ͪ��i��4L�hءdł]�H�*�֡yh*��x{b�|���޾f_L(c�8��5q��3�d�����p����~6�4���S��vF�]��F2�+)�ں�-0Y�Y<H��^��4y������-�}4&!���	�5�q��R�x��h�-���������x�e�"�^�i��0bu��/O�;!p���A߾� &d�����)��
אַ*p�� &�Ό� Z/HA�<U�o��ߥ��]�>��FK�	v;�D�f08���eq��I�K,�O��3��\�eܶST�-L��ȍ�ʧB��'��৭��F�k��.z��<N�'qM��$ULZ?�����;�njũ��S�x��4�=o7�.k&��$��խE�vQ�9`G��B���W��a�=�a��Ǐ䈟�4.�Fa�p����*]!���	|w�:�o����ÅU��X�9k���3F��4�iyC`�q�C�z��Avo�X�NgJ@e�D�������VI�[�'��{�J���2B��+{S��>��Ѣ�ٙ;�0�Ar��Z�A��RL�%�G27��z$���}�[������~#r$�-G�^�+�q��ۜ�S�Jc�q�0�DP�vZh�p�\��۱�w�6���n��W?�QٿP^=n�T��e�Y��R�F:�4��H�\��3����	�!a��4H.�+*[n�������#F��d���"w9�7�vR�d��4|6 �lMP�Wÿg�o�M*n�W���a��}E�(�Hd��\������*�w�ǌ>�'8�mVv�b�����\�sՇ�hۍ��N:)�b���$f��N�w�C�J���aW�I���_K}KҝDAr���p��o�iu�j��
m2���3V��w�n�=��3-���PT���f�¯��e��
 ���~�%̗��{�m�n� �N��=زR�����3�n� �5���M�;BFƝ����vT�<;*��eRܢ�����v-5�u%�����OGy1A΃���'�\|�njs�!������O���N���=?�G��'R���v�ݨo-8��D8�WK�m��$�M^��q��=��0��I���g�j4[s��2h:��j�-�A�E��)���0��=�t7v�KT�n�N�I�~]��s5G[#�i��t&�������ls�$��c-���N�~vo���h �dp�U��>IKOC"?|�����PAR���AB�-�+�8�yt磌�
U�UB��D�aR��#�����Wa�8:�~�X��H���y� ���<0��|t���Hc'��My�8>��/_�kv��캙�/9��T���
DDR�U��m�%�_�"��/�n�̰O w;Fg� L��-�ĭL˞� U�㯽����o57���c�$�T9�W�T�
b^f�P���}#(�ʽ�N5�?�Ʊi�U����X��`�|�����i���$֑e�%����w�%�̄�
o�:��}���YU���i���f�
�6ŋ?;�=�$���t��^��g�����t��P09�}�nct޲�f�}Հ[&�&mv��U���<��^]!��g�0���D:�;�xW��y�X�K�0�����t��dV�B<_3k�1O�A�'X=�������6�00���V��Ё�M������
1�?J�{ߠ_M�^����0��yG��{��!N�7�����IYTϛ��7���@G�^ݠ�G^{�cR�!kw=��6W�*�~�����Ӈ:�
�;o�d��KO��j��*���bp|D�8:lE�4y��I�;.o%U�F�Ѯ#��ơ�?#ēD����_?g���TQ}b�F-)䮖l�~�ɇ���;v,��Ȯ�0ç&�F�ղ��	�����J8��F�} �=���6��_��|E+C;ע�қ<`���[ĸ�"��i�Љ.X���C�:���h>��T)TAWx�����+V���]�eI#��+'*c��+��5j���b��m�c@�Z�<��V����k�[y���^��=��!�%r�,z�)D.�j�ڇ5/j���B�j�^�L����$�v���{�oԮ��v^J�~Ń���[G��ͺ�߷�'2����\1c�R�˥�s$����*-I|��wN�϶��\�H��$�s<���z��l�G�r��e��V����j �|_?����zJ�0�f~�z�&���鮝�F	���'���G�N�So�V�B9e����6�̎ڊb=$�*D��Mr	���}Lh�g��91�̆Z�X8�W���?����B-��tb�z�#��J���?;�A�)�M�y&�~w��E�c��5uCc�l�N���=������h�s~�c5p����I�3���>R�V�.>�Or� ��/z���R�R$�$��lw"�Gͻ,t,�k���(��j�d�#�nA{WM��8ԕ~�5�[v L��p"d�����\��6��/��K��5��*a##�\	2��룶L<�� 9�	U��u>��Nt�5�-f�5-�)DwYd₽4冷�Y �i���[�H	7o�[V� Ac$O�ãL�v�aZC ��Z�Յ��0|5�?h�NE����aV-��`���V�P��#��d�����)^TX��f��b�a,aZ��b!�����H��8�x���)'�B�vvx���tU���M�8�X�}�����t�KhaΘ,���Ц�*A ��4�@�T��-�MD꧉ufi8<�/��/{}x��]n�[:j��˺qo����}X�w�kY��{��$���� "CCP�;.�׽ro��2/�L�aV�U�'*�_�)v��!|��k�_e�����S�w'�1�7p�~N kT�^ħ��Q�YQ<�]Iz9�����Ԣ�\N����� �l+.��ԛFUު�L�kje'1�a�qgQw�B0�܉�Z3����^]@ԝf[@������&�� 9��6 �sG��qu�u݉<�hG`���x�8�ѳ�'Ը��x��/*���L7c�k�/)K�m�r�>�����8�RB�K�6� ,�4G��:ݝ���$�
���G������}�]�q�����F'��[B���!��-���B�R�]�� _��.�a&�L+mV
;�z1�������p@Mp�W��2�J�т��&��V��B��[����H���>�T3����Ƞ�l������* ���0G��XTP-0�?��#������Ҍ�)���J �����BT33F�'9&��;�ȴRc������⤞�5��j+����u��&tK�=0F �-�'!��]ߧ!�K����	G��n���#DH�B �ܔ��u\K� k�O�"�mZ�ae�vUތ#5��f�_��0;qV1m̞6[Ynu�a}D>G�>��V��x֒��fJM�;S(�\�9��l9I���v��c+�)�j�K��v���?��JbeH������8���@���pc��T����㙕P��i75��4� ���Q�x�rWg�W`q�w�<ǚ��\ �z��;����7��ީW��4#��D�Yu�39��WI>k�}g�,?�y&��|���n�
'nG��g`����3��⇓�v�9����n��R��]��>Ob~ i�@����c�Y��@{.�}��Pjw?�p(^��Nc��$fҮ5�#]�5/��l}ojz�\��I*�Zߢ�!Ce1_H7K�y�睁Cޝ�Kh���@��:��YMF���1�`�]C磩�]�V9��!�Bl�,���Ѕ�q���A-��6s�,��?�>�|gي�i�~�ğ��sMwtՓ/��)���i�VE�\��}҈G�R�4�0]$����c�|De�%����a��m�P}*�4�G�g 3�*��Ň�oN�/)n�R�K��
�\��L�g)q-�W�c�h?vۭ�h^����l��hs�=v��J]�v�Y�sd������Q=UR@./0��@�`�b������	�@X*�.�r��\�F���kz����tH�k�pIMp��b��1���м��>2�!�����1�Tc�s�e�pȣ-� B����Uev7�I~�tJYs�0`:�lR	�]���������g{b0f$�����+��6E�����A�2����`Ҵ���ɓ��D�>$d�c���	|*��ؾ�J,�a�O���E���*��[D��V���e����q1{y#���b?�\���o�
�?*y̵p���F�V��,n�Ԧ\DAI�ˤ�Yd9��J��/#�_¼�X�C�P��Q���?PM�U���4X�y�,٨��o��t|rФ|�kM��2�M���\�%9ц�K�X�"��![:���^��/��/Ύ��e6<�����?[@X��,�5c���������"�?�蜞��^ɳ���"�`�3�	NY�Q&e�Q4Z���'��#+~x�^���t���&���o��j!�0AZ5
�,�N�RKT>����ݘq͌�,��w2�b��e=�� �qH^��`�9�O�['#���}	���c�r�P��_z�bs]�o`���2]����PSS���_�ۉ)N�QV�UtW��޵f�(c�M�%������]�b����6�]M�}yeӄI{��w��q��7#�]�〿����~�d�¦��LH��3N�k���؋O'�2�B��<ٯOnK�N
R_深|��c��Gs�m0���t�xS���.n���練=��A�N�xj�3�:8�{��"xjg\�����u]�n�!Gi�JW��H9ǫt��R�bp�k�̷2�|0�7u���+�KE���Գy�A��G���(K�7����ӑ}�
�Եo ��bP�	�qp���;�W��9h㻯ez���_u*��j#��d��C�g��Uղ�d6Z#�%��7�7���p�2"̄)\�%3׏��nK$�+9®4XK?Z�\��aA��\�q�=�sX��#=U7K��-(�a���ѡ�70e�D�N*L�|���☏�5�i���9�0�۔��:p��;�0�ƅ���كU��X{����t߷gA��ب`��XU���"~y�-;�j?� C��$�u¤ڝ�e�m�{��i��5q��<��>Պ��:X�l���cz��Uy(�Z�s�4]��L6G�b�]�r�2���DJ��U��t��5�p���$��_�R��R:��xN�D�����{ ��{�2$��CF����h��$A)��� �[�����+�kN��2fH����kҋm>� ;�>Wwl!^G��\��s�w]����x5^�0��a���L!fr���[Q(T@���븼c6�T[ 2���� ��*)��<6m'�J0&>)��o"L|n>�s��dAZ�G���2�4ˋ��}7�uӳ�F��W��F�,�����0�Hn뀂-� ]�BO��f��]�C�Ś+N���𬒔���)w���p�Z� ;�,�$�%ޙiV���VµjjƆ���T�����6�}c��eΏJl�)�Ӭ���G�B���eH��m��Pr����4�L5\ļbDV/��.`�����T�+�]��\���{p��7��5�5�hv<`D�qh��y�b����O�������O��1T@Ӳ��h+ڳ�tF=,Jh튵	����Z�z���^��ԛ��MwZU���$D=���{���
�����Y�G��y�r;����P�O~܇p���)����[y^)'������/�<���B���n�=����z�Oկ�?v�N]"[�(NGּ��[�,L'��9��B�
���M$��G��+��Z� (o��0�d�7^@�W�Ĺ���D�ԓ.߭����{Áp�W���\��&���h�E��q�~O�@�d}q��8F����& �b{0�ˇ��ڄ�$*��ԯ[�Gx����20� n�����|�'�t!D�q����q � ��-�����b��@�����쏉�ȸ�|���#�rP�4m��tي9�_�	.�8�Vt���N��]'U1��Y��p���8^U��^ϰ|�6֪�i�r���Sm�y�lyx�<�(��IH'#L�5z�<�������F�i�+��LA��CXKF�
?l����nU��Q�B��7� �v ��:�H�g��va�ZݽS�\����hƬ�s��]vz'O�t���q~��a'�=M�M�G�P,+���l�Hz_�5%�z��+�l�͕}s�T}�۰�����>����x���
����y�N���L٣����|{�t6q@�F.���s�ORkk�b�m�͛���t=s��nF��"�SWUm8�]�βQ�eV��9E7Lm�?"&D�okg\1�b��߽q���?t9����z�p �5���N�O�Y7]d�T9����8�����W��r/����~��;���̗Ib��rZ�H�!E��c-MR���G��s�)��X麐��J/���r��3!�z$JU�ܩ��H	Ԩ@tb��tA�~M���8f�k��1R\���~�]�Tu7&�@]�n��c�`$lzI����L# �l�F��C���y�r�*�����\�,	pD��T|�lZ��z��aJzj�c���	ʾ]ZE�Y@$�=$���KY���E6d&;�Ӛ��ȝ<��z�������3e�����F��6)WV�F���h�
����!��zk��fMH�V! �����@�WQĭ�7��	��Nku|)�}D�o9P�ћ�Kt��[��샀i{��i9ޘIx><�`� I K@,(P�z<*;���Vk�g��n0�7 �ܶ��:�V��ă({�CV�xNaY���+�S^�Lp@�lC�|O9��1ۼbz"!�z���P��]d�L�Q"?�J�MJP��ޏ���
T��f��Gc;�p[m�䨓�E5[!�D�6���-Z�u&#q��	�)��:�oW�d"���kG�pF�R������48���}$���.Q�E��Qk�L� ?���]E�Nf��N>�7iG��+E�c�	��c��9σ��~g���i���:7�2�8g3��wܘ����JN����2!��=��u�	�cY�d�J( bUv�KK@�&2���cc��xwxu1'?�מ夽$�W���c��6".���կͪ`W�C>[Z}/"�Ȍrn��r��{���xFHF�����������ű{"�8�\Z�P� ��v���oi����r ��q#�|Bel蟛�렯C�;Y�Ŵ��x����6	��ݡ�M=#��Y��Gw��^��FG�P)���h�)�@ja��a���&�N�'�p'Bu���S��|�M5S�\2��n�%� l�[���]�V��^��?��S�ܴXD��L�]S�^����g+q_'�;���<D%a�)�2�|c�����-@0�U�2��?E:�O(n뷺���<ZR�������R�5>�X��Z3���}7���m�4�Yp�(o�Va=Eي���4f-Hk	�ߦH ��"I�m��;��m�P:������u��U&g�4�Ͷ���%����+���˾mf��Se��~q���)u��6�c�]�_���h�f7���-mQ�������jyG�Yz�O��
}�*6�k��YY��*=I�"[��!���5����2����mu�,br�LGEH��Px"�r6�ίT����
�]�ҽI?�V�|���̫n�r(�J��J���^id8��� !P�I�C3�jlU�o�9i΍[�xH2:�P�Ra`�`�j�� �`�) ����7=��
tm��U	�߭y�E��6�����0Z�i&4c꺌HE�'Ӯ���b�����Y�B�'�4�h�aA9x\�ȏ�P	l�uY�/�0�P9�{4����z*g�ܷ��h�ȞM�F�ԡl�L�$Z��`y��Gqu�M]G�LB���@��Γq[�9J��#�bDCi�0����ږz�u�/2r�c�˓�o�Buj�y��=qC�!����e;��!|xv2��2�[2��-η��P�ixC09�?W��~�B�i��9'�	���|�ō�`r��c�_�F�g�
J�5�r��c
�o�B����z~�SK��Zu��ub���!jXQL�6V|�Wȝ��]�ꏑ�t�"��Q1�̐8��͵���5[^����1�F:�4����ى�m�"jR=UQe�r��
&N?��bb�)#Wư���[��{��+���k�����%'����}*�n�d�\k��8^:���ř��57MW^��gJYC��`��~�y�����g�ӳ�: =m�vܣ����11&�~�ISćU���G�}�vC7n�;�c��^�L"/���̏ۚH@j��	��s����7�jn4�;A�;�K��VnT&�Ƴ�K@�R�!-S	իxe�Yr:D'�M��~E��5�d�G�D�wF�;��ngnYH�Ӽ��Pǻ�D>b��!z�ʋ��d��%);IM����'K���Ni i�B���3����!��F�;�?m����71�:�* Њ�c6*�a���vlFNFA��%��џ"Ģ9c�(Pi��A=�Ov���/�蒩����w���̣)��i�7��� �u9��utX�W����n��}qp�%���x㤐(\/Ј��A��-C �m9eV������\��D�6vjp�Hxfy�Jed��g���-.��iU�Y���^@�g2�E�N��s�p��X�K����uy�4��֭b�y���#sX�9�d<q`�"�,	$�	{e�rqgH�v�Э	g>������W(�O��zU����4�ZU�JNY�L�F"���.�<��Y����VEwsx2� � ��V�;����bn����D��@W�p<=o�҆.�"'����(�&���I���� ?���]���p�y��<'�S�e�d�_C6dR�t��=X�@,U7��s�*��w��9����Z����>��;������ֿ=�� ʞMz'Ic��S�rY ��/�禞}���>�%����tmD��,�U�v���G5b�]xj�3��n������p�'��T�e�a����+X�G"��
����_����:S�/ñRo��%'{dg��u��-vo���-���dbE࿆@�by���kus��1W�ΨT1a�]�	� �B����4J�m}���_�����;L�m���F.��M�"�GT/Ћ 3��9�p'՗��ƫ�9�Q ��ۑ҅�Mc�4�H����AD��u���:���O��������@��u��7�Pp�A*������{��UCɑuO�
�'�m���'������LYDR�Sz��˂GY"+�b~X�p�0K�Ӯ�ƚ�h4s�&�fΎ��bI�F�p7�~I�+��n(nb5�0ng�}��`gYP��nFsc��tU��!�؏����va���N��<?��!ܸ��c��֟ox0�~�������?����t�r���w!O���eJ\n�����'�ޫ�˘-Dff��;=�:�[-�����8�vv�c���5�k������ �ػ��"z�RUz�{�"��ßQ���22F��ߋ?"ܓ�9�cӡ�9ϯ�kġ��1�cJ�B�� ��5I�5-�ؒ�5�Ie$��v��h�}�~]]�$��vu��M��v�{��l&����3�]#���G�eKw�/s�v
\c��|��h�Y+��*V���n+T���'Fa(i=��2���2N�P��֠{-�yx~d��;��A������թa�W.'��n�>��h���8G���A�4��s��һ_��g*
R�-��|�v���B�4]%���6����#�1��L��ԭ�(���+������D>3X����M�(<��K�
%V����Rrq��WC��"�a�����Ti5��}�FB=���x�!�j//U�#�գɲ��ȯ�l��z���p�ɭ}HE����s�忍LM^u�����_zW�R�7��$e�[OgZswVyI>�r,�E��`�X�҅��Y.�K�Z-F�N����y8�,�7Й०�Z�!�8Vad	���t��7TI�m���k{36����Գ�I�2B�U6�̷�����l����"&���hd��P�z���bӞYW9G�1�K~]�.��L*��D��0o�_/.O�ɄY7̊�)Ys�DRos��c��M�M��nt!ǪV�M�v�[���G-)�E��:����
�t�5����O6��D#�>��ٰ�����2�F<��̉l*�͋�{�R��%�����h%�~*cc=^���pπ���w�݄vQc���݄���A�_��'����d�^���Ɖw�`Sj��0�A/��V�,�Є=8��)���۷�,|�`�KZ�3�o5��X@y������uC����n�+l���OKI2!���q�}����|�X�a�b�)hۭ��5u�`�ja����E3�C�z[������e��h�!�վx��:՛�C�&��X�"]���� A􉰑�6�V�:�F���^SU����	�s�Q��#me�\�PJt�?Ir웙��J���,��r6}��w��>Ǣ��]��@�Ī�OŸm��V���8�fľ�0m��x5`.�Fk�7�>���'��y�g:̶H���N�Q&����?����9��^�26n>�bt}/�3�x�Pn�<����k���XNX�0�-?;��= w9ɩ��� ��ܘ��F�ț]~3@[���`� ��)���n9�>�����g(.���V�׉9�u
q��̕R]t݄���<J�I�ߴ�R͝J{	��q�[�nZ	��S�o�D�N���@֊ic���"2**��Q f��x��1ǟ��E�j %���r�6�Uh��Xh�G�b���=	�����1o�7w�a5a��;�O寻�y,�O��E����E������r�(..��{<���s߅�ݓG��Ϭ8pA̅c>+�!PˎPd�Ŕ�rK)���e�O+��6�>\��`m[�����WJ�n5r��\A#��q�tǸ蛾-P��KN��PhV\' 5ݑ���{�T?��"�v���Q>��E�z�|.��Y�d5i�����������y�h���	�s,&�*��@���&���9L��G�������}~��w����f��p��7�
�&�*S�e g	�h�^	ި=o���а�:�^;�V�Z��6����"����(��w�����C�?��d��K'�&�.�<���f���Xn�6��!P@�i�p����.y�����r��o���>S�<�
.~V���~��;��
��y�fN!�q/-��3,%��
���v�婘�������I8���M��Q�o,�Ɠ��轂�L�[���ҥF!�����{n��
��C��Lk�=�Ϥ���b�:��ls[\n�V��V>���je�KIρߵ����Qi����ON����+�,��H�)�ئkēw��x�B�_�h���)��҅f	 {K�UZ\3�gݢ�U�4�<��ё��ί:F�֖��d�e-������3�-�(9�t���m�b�B'YV �Ow������C�$�ӣv���3�*^��u' �,�ަ㗴�3�:z�^�1�S���|D��?�7��}9�-�d۷��]h�b^�v��k�ngs34w<��o�k%r��1R�A�䁘
�d}�p���������\�&�����6-玌�2��X�B���A���Oa$�v���Y�uE:�Q��!�&ŉ��z�/�tX:?�b�L&�k��a�~���d��Һ����n?(J��S�����
 �*e��G�?
&RJ�K��T}d��k��$�����2��\k��p�ra�4�e52h)����ݕ��g��߳'_�q�j�|0})yMUח�>5#5U��D���׉ۊ�k�g�ӝF�8-�a��ڊdi��m7}�Z�D&�#*�O�ף���[kPZݕ	!3@��:���<N�$����"����fnՁ��r�0��ڻ�˶�
R����*��e��K�U���6��YQ����y�ߟ�'9�'��=dT�IVueED/�K��lS`��l��o��z�i}�")��=p�	�9�]j�/x)��A��u���C�
�.ss��T��с]�� _��Pg���u�x	�9�s���0��"����	&7�)?;��$!��z�N��<��B�ҟ�P��1� �=d{��YU�P�hc�,��yiLt{d�b4��3@�9�>mPo^)o��d�Ȉs�L2���]�\�������7g���+'>t�{G3n����GD�:�s������i����nf]B5x�J	�;��X.LU��vt����G�ueI8L�����6��J�:��g��w��U6�ۣd�f�V�-��{��MDE�6�p�d�}+�� 2U��$4�~�'���vb�B)m��������.hA�B@�O��-9&Q�~�� ��%Ji4�p����P������Dw<�����];v�IK�7�����Қ�8��3ը^�Ǜ����y���9��a=/|�sP�|�j�r	Bo-o���ɔ�l����q��}ɵ ���ق���m=7��+E�g�a��U�� ������I�\�M���F����tt�R=S(r�է�C	P�̆��"<C}H<���
3�$�]��ܰ�_w�gi.�� ����8���{0���B�r����W�u6'}���:�ml3u�T�
�I���[���#v��� wt���~2�J�G��!�6RI��ُ�j�?��_B���	����Qs�P�m}vY*��b+�Gl��#�M�$���Iq�{`%m$���LqA����6�α�R0�����$X�dp�M6{;�7��0@;��IW+M19��@*�������|��=M�:R��, ��	"�K��_Uo8"}����+|7o������B)��3\��S��vD
���z����5g�(1�)��;��"�6��篙6��b�W4����N���z�f�V �Iҍ^=�0��+��Y�ˣ�>�vې>]�C8�b���0`����??��(�qN��	!�˗�ȝ��vr���NP��H:�)�	�LWW�cHi�Q�@@�m�O�M?�Z��;ؼ,^%���z��ϫ4ȵ�+[��Q�4NrtO ;RgO� �B�Йj�8��)�SՊ����n��~.��JB�-`q.z����U�M;�B�o���^��|��Ȇ�9��L��WW0IJ��(&\$`?��w�r���SN�����M0ߥ��Ts��P�)[5n�i	%@{ʚ}[\���[�'g�y�[yMbfl|�xi"*MtI/���&��8��E~��O�%�mൊ��r�� �/;F#*QrgR�./��E����x^T��	��EA%^⛣��)����?n,6w\I�g��S���rP��]��|�j���H��$C'LR��>'�T\/5�_�l���x�J��D�Q��ʰMu���	�X�H�J����9B�T�^��C����Ü޴��O��n%��AY����HC�G!�)����s4FHn��P){��'2le��)x`x4;���x2׭T�S{�Eҋ��'�{�^BS�
�*�n��M���:�޸)����l#��_���~D�:�%� ,�oVB]�<%A膉˟}��t/.߾8z�V3mL���SV�5�Δ�kȬ��b�>�J�:�9�hǞlb��{������'���e��ҬO�w�r٤�Vɑ�#�{�UGt��̋�>#��y�|��P>�����z����ӷ�� �'!_�V����i��Q�>l�Qh�\�F�'$�UtT��?��̟���M�x'eN�A�(N>���6���	����72wj��'H@��A�
0�4,����×�0�)�7��{�$v��S=�(,�@e=�?�Ւ��Io�6	�hK[S�{��)�\qw�ג��ʻb��(�c��U���f��5�������~3�<@	"ػ�¾���;��J$8U��z@Ct��:'� A�vlf�L�z�;$�5H�Ch	�o��H�� ��c��{��W�q=}=�a�h��-=��N�E�]ِ���&��w���h�?�A+~q%�vس@<73n�abf;�H1
4Y��>��m��L;Ed�n��"�k����di.���V�e��1憌�u#�G��O�2��5��Ë��uz��ْ�׌����g�A]S]*W�EUYz��~}��l�ֳ7.%}�1��k��{��(VZ٠@���}�����U�t+֏�g?��]��ߍ�5Ex�8�Ѣa�战{hWW�۹�Se���k|ZO��n��9s�v9I_f��?b꨿$^�;Q7���iL�P� ��.+�5)��H='q2�X'��L���wO(D�����Q�3�&�
tN�y�%o���rajW�L�=� �B/v�#Ki&�w]��*i�j�{����}W�J��уj_\�"i;)ނOj�����'ܢ=�'��RKƾG�����k�&|�nc�A��D�_��1+�q�y{�=69H�<���q���`�K�h��2E�-㺀����W)�B�2�Eqm� ⛹�2|P<'S=�z��B�*��)�fѺp�3�k�J���H����ߐμ0
��h{"(:)���-_��6y �U�8�eB9
���0��}�r�A��˃�eM��a}�����q�6λs�Ƚ(�>���[ݐ�OaGTG2M����ҳ3a�|0��3$�'??�������mz�>�	]>�0�D7��6�j�������h�"���B�^���4o�\����/���!}^�A�����2�Q��Ĭ�*l�j��am0'��E%?BetД���m®
��X�C���0�Nm@�E��2F�m�`��A��L?��r���	�G`��- #���-.H���0�'{(w?����$���[Y9�0^*��2�4�������١5��G�h��}=ݳJ�7VH�� {D�d%7P��	�OhT�ϛ��1ޝ!_}�	�~g�ot�o��l�xpN�&��Zzd0�.⯕�5V8�[ٶE�~����H��S^��0��SL��ٙ�z�C� ��uF29�[������M.RO",��\��7�*"	��@��SB]OѼ �3��Q@R��}�ˮDb���e�!7\A��G⏍$1��k��,�, �l� 3đ�[�_��!�����FN���i�� HhM~��״�����0�#F� ���Q�E9��z�>�����=ha�J�����)FT�Ǫ	�O���Ē�}��D��l|l���P�f�ľ�����e8V���# �6�@���dG�!�Ξ3���x"HHW3	旅����T�-X���Ҹ9^V�G=x�j�-8����\ Q����d���ei����W^�F>�$r�*�\��	��y�QEI�e	���f05�ۙj��Uщ��Ha�z!��G^m����J/�4�t(H���k�4��++�a�쵚	3%�
��0R��g�=���ӯ��K���:_�Ay�
ȃ.TԒ��T����ަ����(!�2�6ˌweq�"t��k+��؍��Z��	��QD�'��t��LJV��F���<66��5���E��Ǟ� ?�!���)ߕ�@���*�J�h�®�ٍ8s¾w������E6�Y'��a�U� ]���I��PR�o�"��*�jhCͰs�0�U�oy"����rd[�{Oyv��o��C1�
�Hzj��-�U'`3�E�v;OQC��	�(�eaeie�lJ<V��^��������c|B��9���A�|`ɀ3,/��G�.�v.��gx����kO���Ciˀ}�$�WN-蒺�N�M���3���(嗰��i�<����i�ڿ�Id�j���ISu���P�����+a�@Bu�47d�4��z�f��_�c��O��1�R1s7�8}x"k�6����>6&����Y���-G��X�u�#��b�p�Z'ω�w��VݪAN\':�1NZ4����&�N_K��6�g8<������<�d���f��?P� '�wʡ�8�i!����^��ܱ�P :N*��P�����-]A���g�������^)�g�f1Ԝ�97�Ё�G(�v��C���B����[�S���F�A�*�89�Ù����{����SxV9.1V���` �Z��Y���\B�znj�z�^���A��yH����B�r����L2�m���|��S|N}��Y�d:Z�xm)4#E2�qiF�8c�j�F������`m�+�Q�p�&Xs3�@��$<jW���;��9�W-�ó�P�~�c�:р��	���̳�"��Z���Ñđ����3q, ��&Yܙ��΍�<d����iJś��+��ޤ�MdЯ�c��kN D��M�m��Q`ʳ�S�2�cg�,��5�;]�F���;���7�[l����T%N�Qq���'Q]��  �0vK=o�*��CJ�x���+�0���*(���@�m��b_�1p����;�6F�_�OK]����"Y��?5�z6��\�3 ��U
����eM�$I�A,�9SD�Y�P�>�����E>y�f~������?�k/t~�}P61ܕ\�/��h�{��%a
?-�Ɉ�b���0O�}-��=<J3��d�
�M(��1{� MD�}�nR:����5Ӓv�E��N�A�� ��uy��1M_�(E�G�l�[�3;�ё��:�������'��g��O������4��D��l�|`ʴ>0����^�U�B)Q+X/����j�v�KHu6{C��ա	k��(�	MV
äJy��%���!�;y��,�:�5CZT9�D�>�nY�n�|G��9��GZ��D���"��3;�W�W)8�Qw--�_ B�66'�~C!Z
5h��͢>�V+^io{�cI�{_p�13��	�|Y��%� �K��!����h�����[�; z��Ƌ�n�� T�Y��LZ�s� 0��H��ð~'o�z�I
��W� ����W�E��m�뒮;5�G��a��U"e�,�@�Q#�Z�u�{.�%~�M��V0n�u�j�����t��3C�&�sŜ4�&{�<��@�;*�Ѥ�b��^+�f�?Y�$ސ1de-zt)�7�����B[$S����1��f����Υ�Gnwv_W�ּ&���EZ\3L}���05�nᑷ�Gw�*S��@N)5X�,�a'c�t~��LxaX�q�x�5��=g'�
U;Hۅ'Y��Ȧ=� �B4e�pj�|�뗵�l���5�5T��g�\�F�gEfO�wC�	+Wkq�j��6�~��@� C�^F�(�� �i����cس`��m2��a��@�H�賖�٠v��ɰ�8��`e�e���ȩ�1-�0�.�g7�6d��O�>nQIQؗ<��w�������L�{�Z�[V.�ci�镽z��DD|�EM6�����D ��j��1���iu�-���	w96鷖r��r�f�!cn�RsVik�~��pd�sB�`0�����{ǚE��}�}��@��]2��L������/��fNM�q�:i����Q.��1���2�z�@���QS%�l���j�ֵ£c����ɴ⢢ڞ�b���>G�S#2��\<�H���J��,�ä�J����r,;��6+�7%��n�)X�D@�5�{��N�:o%�z�\v3*�2�F�YOݜ�g�X�*.}/�J�1�a!@��c�X�m3.O��"H-k~d��g?aRB0c��h��׬_���(����_��P[0���J'�:J~��\���?�a`s�zN�b��-��<�R�����7�ݕ�,b�>��}���ݘ��g��wz� �b����X%/ҧ�}�a.<2p]�!��ĩ�ֹF�C�&+L�LW�*�V"���`�T�
,bӪ����'(Nw�D*��l�nB��`P�n��;�	/�TXN`e����ኄ�<8*0�߀E?ɓ���*�B�
Fa���4�U��w�d>�֒��l�i��o ��Pt�p[�X�t��w��Th'Orl�3�PJ���r�ʧmѓ_�,�B<���w�Q�m[��_��(�I'!GMٰ8*�V�,cc����V��#/8?\���G��?��?8@q�z6[��P~;�|�����x�R���כj�����O�Nֵ:D5�שaG	���.C7�B�/�j���m��M�1	��k�P.xQ�̕��W���=ߒ���>������Ӈ;r4ȃ y�=]?�G�h8��]�L+��fC��aeg̲T4�e�"7\O`e�Xd�?u]���q�)\�����}�&,���rx�F��}��B�0�*��A�.m{	�E�y挶���78f��e�ÎU��l�jq� �$h=�s��Y؂_7��i�쟦~�p~)B1���Bȇc9'�"��ĥ��յw�sy�MԴ���]<��I�)��{��V��n�|���^=e�M�c�דy�#�lLQi�i2q�i�p�: s�=<������w�
vS�`������B����XJ�������S�>�.h�yF�p=1�ʄ6�%�>2Łi��9��N�+�=&��"��M�c_��j��ڻI ���63�����!��_��յ��#ݲh{���ȓ�jNҧ1!-�4���P�,((O�ϕF��hy�,V�('��M�#���+�ȽH�pOք
(��N`KzB6�a!��ªt>>�]͟�܌�s��#J���d��4���[:�ǣpG�=�+�#���^��nG>�9z��/��J$rU�Q^g����lE}+�8�˲c�i,Ԯ�����+�I>Q&���ԳH|;S�u�I�z�q��f��7V9�r^�w���P-mC=@��W��R�� =l,H-�$߮�Cu�f�6~`�~f����!��d% |B��ȺN�'z����rtZ7I�P�.�9�&̘I�����O�j���?�۽�[�,��Q�r��/����Y�;$J#�\���?j��`J]����#;�E|ˈ���3=��59�Wnt�
�^1!���%�����G���[ʫ���g���8/{}�n	�V���aL�Jla� �Q����o�?\}�=�_�͸�B�����n�`�Ŝj�9�N˃�����%^�wi��L�2���[�ۗEJd����Z�k��5�IH�/���(.O�}Һ)��W"��+P�y����p�gR�'q'+��IsR⛷ؓ6��B�+�7f3�D S�� �e4p�Z�M������E���"���۹d�pR����ة�z�_�9t��삿��W�(P��BA]�L"�X�е��� =��=o2"��nN��]�$�'�6�d�P� �~ �C���M[������C-����T�
��*��p[�"+)sTd% L7K��T��T��~v,�xЛ�uj���lY4b7������g�#I�lq�܎DG�'G���S�	<O�&pH�#��_ȺQ�gx� ��1�(��j�j�̡�.��g8g$p.��΄��O9���)����Я���V�G��N� �����#�湩� ��
��N�(���t���-q��ʿg8˦�D���ѡ��ئ�YySȮ�R�#���+T�i��O�d0S_@z0��$�z0�b\;D���>�𐗎�&es�eʌ�_C�~o�X�Q��sDa�8���Ru8"���#؞=�B��-��i]{���i�=�[ ���d~��2A�N����x�A�����^���A^wF��Vv����]�Y}�����fNɫi��u;��G��U|k,U�Nb��iO�S=r$��z�.@+L`^�F�/�UYn}.�*s����v��n#)�4�F�L�&3�<P�N>��C׵�	����[@��q���;��ݟ����ɋ)�H�.y�2�>9=�B̷����j	A7�SQ�ۿ�F�3�E�K��C_,,0�̍����o��p��L�Vh�N�����^���g�`�q�.�PȎ�liq%ڑ���1�J
l�}��i��_o)��,ړ��mWƒ_��!��¦��3E��t;jo~�>#�̮oC���a�.�rXԬ��kVF��b��;P�Ysg7&�D�w�u�/�����to�׉i�}�vC_4�����Ԋq�r�_���?���f���џ���*Q���P|�j�$R�ds7�UQC�,	�gK�
�fl8�o�� ��$h��AkU��vKDS����e��q}���l�C_�a��[�@�]5MenjLΫϏ�n�N�a�����ha�C�N*n#8M�X�
5]m��K����"��Y�9�ó���=\�A���rG�-B<��k��Fc�Z�<[��B��`dG������fv����)~rs�!i����l�&�AC^S����tfB���f6���q��'�<�f�DM12�5�iS,���ߜ�f�P30��<e�ZB��	Ǆ��3v=A��
/=�>4
Ф?�������z�tb���C�u׸p?�o���˚Ij��Q��B7RsO�-+��U쑥亁'\J^\S�g�=�k_���>��ԭ�9�K�S���4�0E���9 C�5p\Ahؙ��B�b3Y�k�	�q*�?yp���K�X���sL2�/�����_��4*vx�hK+!H]�˛xxI4�Z�DZ_�\��3þK���������4�(8μ��.򟈅���;��-��8,��ظȕ��[{8�qV�mlDp�)� ӁչG�M������@��=���H��2��kM�)�Yx�Q�l`Q�U�@1�""~k�X�p�h�򌭉a.��^1�3��O��"炗����7�����jyH�I�N.3�Җ�hb<Jg�ƹI�k#�c��HI E�\��g��z�ɞe����ܺbR�ɹ���q<��gň�G	�>N��6��XYY��A	�&'������$xt��<M�0�I�cۤQ/�e��$#�Ȗ%6��h��6��9��P �.o�+K|	4�,(a��Vu�B<��K�	�!�Z!ڲ�Q�
"ڻ̿Dl��(k�,.V�������ϴ��?RbPy��{������9��U�z!������A����x�nG/� `vxH��]}��)�������&&�m�P��t�!<﨎v��t񒐯�0��X4xE'��!�T��xPcU��w�mN�#m�VOט;6C,�kx7����Q����6�!w*�����1˃��gsgT3�F�<���Q$���Mw>�B]�dAW�����)=<�Ab�f�Pu�q���k^+w�c�.������Ȱ}N����ͯ��`��^��uw��0 ]GC$�~zaJV�`ʾHQ����t��e�P�J^z��Β���=@9������
���ˉ�+L����l ��XaG�]�K��֟��b��J��ƥ,����VV��όl�*q��i�ǚ(��F������׽������5~��&�UZ��l�����u�L����Z�7]0�Z�Q��M�B������_h�6���nXO��sG��Z&'��;� �UQ���d��}"���l`�W��d�Ğt�¶:p���}?ϊvq�81fɍ�vl����l�U�H�0��$�V�F�4ģG��tBr"
ʨ��/*�)�Z��T�U�#���w"y�3�B���[s����s��p��X���'�"�=��k*iL���9s���ĕ��-w:��.�2�@þ`��y��Д{��j)�8�LF����I��M�%���G'!@�瑊��m��c�4���Fw�g�c	�}$X�C�.�sT<]G�D�S������q�N�6��S�;%<��K}� ��g���V����ehy�B�����Ƚ�Lfbu����lc��z��TUcE��L��,A�8/(?���#�ʖc���Dv_Yxl2�Z��j.to�eف�]���t���.�]������C�ȡ�~��fe{�U���}ڜ���wq�Z���:ה<�3wIk��m��,m���%�e��F�L{�Ͻ:��>�a+61N*�FnSq���-������*�)���4J��ܣcܦg��<k(�9h��j�9ܽ�k!$@ř��+p/��4��B0T��Gd���CO.b�ԕ<�a�{�w5�CnVɹ�Ww���M��]�CW���Ŷ���g|��o�|0=�.E��8�2���(*��?Vf]����t>���,��]�O� N�%(Q
�&�F�!��gЭ1]&�)��/^��-0�3��r�qe#Ꮵ���OQ�\g���/� �s�0����^�(��ɱZ�EP=����8
��x+��n'WU�iu�v)�
;�?�q���Ĳ���,��s�Ȭ����aOH=�HTg
�!��jN������dvg�m ��Ci� �� �Bp�ʗ���b�4R� �u�m�vf���UԻ[; ��@^F�m�Q����Z��
�k����u�_�Q�l�S4xk�{#ht��9�9x���' 8}M�}��` +W��G�O6FS�TQ�G#����Kޚ�y]�[/M�rH�u����u�	t����	�#�@_�T��h��C�tנ�⤳���9-�O�jOy �A�*�B�UƆ����#^U-�g��@�X{Ξ������ �<�	��]ש��#q���Y��Da��Ώ���g0�� ������~�����$#,#����v5��7�؉sn\�m@�u��1HLϒ�tn}�^��m�R��}�� p9*;�P�L,�+�e��m��&/h	S�V�#`���o�ԎYD�b)6�}�r*�0�*}<��U؈��C1�H��_�g�,��k�V���V�5�cVѥ����&�x~��֐�S����)�f=���%���1.?W��s�'
��+�3d���YE�Xk���0&Ёk�Y�N�d�����^��B����ʹ3��Qe���|��B�(T�`Я�&��M�6�R����Ԛ
^z�a	����?�!���y>q�	mDr��]"Ic?����O�F1��y��m��(�o2�xg*�N���f�8�-��
���a�	�d��;Aܲ���K��F1��+��3��1]ת�-<���J��a���b�L9Q���r��t������r_>_$��E�eoX�*l@`���&XB.��E�0W���U��w���d�)�E`9-.ܳS&�i�
AiS{1�Xܰw��m��F2���_��}�=��)�L���;�����Zk]�Q���R�l���7E5�K8*Lv�����8V�g�����z�Usi�^��=:�Cn�$%�S�f�>�hj���]X�w�ʰ}��#zYE��f]�X���	�1�Qn^IB��md���4#@5���u=5r�y�')�y����m�z�Fg�Ί�ʦ�W�եO�D#����V�܅�CqP~�2})�T͵��Mn�)�a����ݖ"����匰�dP�Z�;c`Xt��;��n�	�Q�?z�0�R���L���<�K��9���}�bt���BUO!5#�C�4��3����A[Q����ؚ�pv�XR�!G�c�H�n�����:�ȎQ��J��ᦏ4�������d״�/�B�1���I��
���0FjcY�+S_���E�x1�`��˯�g���ϣ�$I6�	c����Eu�AT��5�t�e�s�?���U[��^b���BVh /`�X!wn�[ψ��y��f�Ψc��;�Jhj%j�K3��*��0DTE����k���żEY�Me�ħ��_�C�,��v�K�]5e������f��d�w�T���ϑUԷ8ѵ"�.xq2{�Ƃx���,�:����	����7�:S�d���b��~5����� P��¢b��
IJNl L�┱��%@2|K[�b��҂�E���a����A�M�T�*	��%��}\����)��</)!�BJm�f�-�����Z���~�@Pl��i-%D��2v9-�X���؎��+e$#N�S��Qj�G�@B��:<$�{S��u0	����:�'D.fv� �0C��dB�~�p%3�6���� ��#[�B4�5LY������>ӡ����rٓO�+v��!�������뮹���%�U��%�����zj�b�t�����?�j��U�������E}��hVS�>��ު�ǿ� �,�Yu�����s����� J���a�yws�ŅMt&�W�g�/��F��v����1M��Q���nX��w]����X����gn!�.�_���!�,���T�O3��w����M��4H�܁���(�C
����[]�D@1��u[�[��eV4��6���Wt�'Y��W��>25����&#=f�CM���^��B�7�ɛ�tP�cf��;D[0OD�����,O̡�h>O�b��P���}������`�������
7O&s����v�|�Ą�������wqG9�q-3���,h���H�7o� )� ouQ�&�Y�_�$`+?v��ip����v�NURt�_�c�2����4�tp|Xo�G��!��bk��%��G�{�G!N�p�p�vh�Ј�n7��ݑi�
5��-v*#SD��`_~��)�����@��@ᭌ�u���jy��5|�m3���_�/�g��G|7q������ڎ2�M*���w���P��@���Rn�:6��"�T�ʑ��,�I�h�x���W��5�9��n��.GW뺒�5"9���]8y%�_�L�y>��q�;vG�i�hX�:+�R�J	������|N�q�;��%Y_�%l���{˫@���F��B����7KT��S�z�V���9s�7[�]��[�,���5fŶ�}�����Y��R�F�н����wEA�����'&���$Cx1H�2G֚:2�Q���C)�ld�.56��e� ��=��w�n����lܺ_� ^kXl�1�� |�-��M��pD#�y�Ȭ�Ġ��B�l�?��������T�s����O����ͪϒ��v�!�~��vl�zN}�1�D0G�	��M�*LfX�����I��������}\n�D�b���a%�6>wq��b�'`��]|p��ϯ����T�_	�a����)�A?�#8$�J1P+�1������1�h��NIϫ�� 	�CA��v�ڍ����2����}��)7=��kt���f����v����e)����ZEk��l^��<=ڭZR���	>8^H�_h�#��<�bC4���/C�R�I�����b��A'T7���yI���^#w�ʼ$��&Z{^Q�(�����?���B�b~be��2�z�u��^س y���#��;*1YeNvW~سJ骟�n���I��	�����흈~@7�]v
�6�k���_�Y��R�܍�oi�-~�V�t��E鯀�\Iڕ����tؾ��V�7Տ!"�i��k~��U�>8������Δ��%�h�����<G*pwcpK�޼���`%��BG����&��ޖ�����)hHlR(g����j9(�ڷ�(�u{� ��T��r��N4WB�M��@��`�2���}�m�pNSc7��,�����`�����>���caj��f2�h���O�@�<o$,_��⬅�_��k�����ǷK���l��Xa�t�Ϯ��I�"��zUeI�W�RU������n��W\fj�j���"s,:o���֨ T��}iLy�O�z|�*r�M�T�Ī���Z�K�|+��>w,�EI��"���!g�{����'�jjW,�J''k��O.�5h�}����dn��;�
��hl� 4z���֫5�b·fG1����ݴ%{}����S5k����Sgv�/�}/ц5�r�U��M�+��k5�F��+C��~)g]591PP�-,.X�㿕�R�d��?.Q�;�
��,_,M�J�+���	���=�����rA�y':��1���ϥ�����DfI��X��"6���1
/}�����K��3;�[\/����/šb#<���72c��ibGF=���i���ä���@��ح�lr�׼�M~��f�_^��r�D�fɏF��/�d��5I>#*�a�s��z�>�2�_p��`w% �{$;�;Խ?a��G�*�j&��bN��%	A�o2m�˚Dj_�*Iɧu���nj]gA��$!�].O@<�}A�V[��A���Z~,��y����P�$a"�C���6~nF�s&(�*�9�v�x9ęAݩ�.p��.֙1�>~J��.ud'�����3<���"�W��2��ZO�����k�4��ж�)L���Q��b��)ٔ�^V%8�z�^~o�<z�3������	���5ʛ�2+Ig�|d���!�Ϗ�6qa���Z�ߎ��B��%:�����e�3�i`J��[�}�`Nյ�4��b1mU�ɦª��R�bdjB��J�3���v��?v���c�M/�G2�j�O�sj|?��R���� Ҏ)\B$z�YJ�PFT}둼�	{Eq�]��;��8P^�`�Q0'm>���Z��"�V�%����9*���n仧ܙ�1	�Dv�^������q]�`B�d1b^��/ �Y� i#D����%����vq�&��<l�<�h�ݵm+{�{oȯ�`�М��v�%��ʬ}�	s�֢�~��M:��8�5�z�,�U)qW�,�] *��ߦs��bB��h�!��tA�ی���B-���}o���0����5���*VÑ�;ʢ?�9�4�����^����P�k=#��ہ�9���&w>��j}WC/tfok���ѼW	c"�ַ@ �����Pο���U8��x�s2ե��{�?D>)M'09�p�v��l�.�ln�m�u'�[/u}�S�`����j����xY�D��o�sU�Z �¿}��	p��O�Y�Ԅ��TׇqG�@�>�����Q�2��O��� ��~D��30Q����	%S����H���.�z������3a��&+%�A����OҬ��&�
i���O5�x\k���v>�S�(>����Q����y�&���$5�����[?L� xy�����q;�<�J���ѐ}����Fl�+0���y@"�C�b�>�o(5�ȉ�|��6�s�vJ�7{�G�q��P�X����k�t��2���l�h:�P#vq�J�+�RR�WfC1�4cSX��½�?�7��f~#-�~��S������4׶����P������`�W,_p�S���qi�Z��I�~���F=���,�lZ1�+���Y�5K�n�HITLo���Lt<+��!yF������\�[�Q��@�
�
_��@��]�p%i��j<qs"
q�zu͐`�������ixi:J�T��/(����~	0�]R��*��L��,��;�4Ak*%Tm�lZ�%��PbbM�"k��W@1cM��z �ܫ��`�LHe����������W�Ŷ�v��-=b�=�74��B��|�����:�m�o_�d'~�t�;i`WS�#�{O��X3��dSx�O�~J���U���25>��[}�K���q`�rFO���7�!�]ʸ�r텩�.O�+!�qE��D�գ�)6�_�XOќ�7����l��aP� ʴ���-�Ю����Sn����2AL>���f�m,�G��_3�d$�Fx��}��W�)�g>y��~��_?H�i��+�P�E��N���9�=4�+���w�֪v�����jx��j�����駦,���.9�v�������d��Q�"��>l�	%������b�E�x�ڨH5S���>c�Z���X"z�רۙ�[ 5Y0����vٺ�
�=m��a�A�j�cIܖ"��z�U�ܫ��޻���`�>��Oz�씂hI�֞�Bo��K�r{�$Y�~��\@.��C/�v[�UL�e�Ox��r�O'�;����R	`�O�}��ͽ����DG׃��k�/1�*TO7��wXw���y�I����T�C�D���wV
eY�O����LP)��%
��C8�0/.��AS�e�S���Wp�Vn'[�!�dN�����)�05�$jX%��8���9^�Ӳ��,aE�����5�#���*��B�̋q:¯#+���js��L���K�q1��~VV[��$�u���t�s�X�I@҄6bˡ�|��uXnǦ�U��{@].5I�����"lzY8(h���2o݃����S`�s&
@�p�	�S�2�;7 �d�vO��s:�3D ��)x-������m��u!l��q�;T��#��m�� ��~��.V�<%׶�ik.��>�z[��,�=�>S�z����k��G���7C��3b��r�))$c�D���ltХɣ���Nf 2�T�͡����s�n9�aYL�.��\�)��(k�o��)��I�]m�s����5��g2Uc�A��V�����b��&]˯��rxJݑ�Z-^����J/�6V�3�h<�5��9�j-�x��)`�����]1��$����9|򤣺��R����ZI掳��ۋ�U�lm#ݻQA��ԃ��;�b�_!�������EnW�Q�zj���c8ߑ ���g�V~gլ��2t������P "�|+��E3J��C��{z�kkRŜg�B:�-�s[2z�v��g�!���_�Ԯ��X9���ig9m}: �1|�����c�M����dv����=��FY�8���$���	P�NĶM~Q�`&{�hJU�)���3��F	�r����5��Ei�׵~��Ԥ��^�eI3�#r�̬mD�O��\]+�IVwMjh�܄�`�5[U��11ʚ�Qym���E@Ðc|nz�^l���~��孁q;w����E���zǼ��_�4yJ����.=��w��A9{Ų��_���#�c�	���P;�����^j�tY�1�#p��֘i5vpZA�˟�G�;�UH�=�,|R����e��ݴkw�Z�L�5xv���[s�{ǏO41�q�ka����T"�V�JZKwT�U/HQ�-� ���7���`���o�E��=��5���^<�H��3lF}�T��X��s����\��8�r���\F��"@"����D�Nm�=0"	� .�R]���]'dro>p{jI\#�T�z��:Ђ0_�%4�Fn���ct��e�4uL�=���>�B�=�6�9���??p��3B��b���(/}y����	���}Y_���2�.v������y]��e��U�-��&��LBg�%�~��@�*4U&�Y��^LF��*�a-��K��+2P!�aў�ީ���q�R����ֆ*5V=��z�l���o�)�װ�H����=g�������C�mPOW�����h<hNqF��
L=�^r�E/����V��|6x�i�qB@���.��vڕ���J��_N�7���! ����_���jt���
�&0Wm��C�0g�[Ѩ���=��h��V�nW�j�����U0�:�|�jFΥ�$|�$�j�=�'���[(�~	2�w L���" $"�]��Sz�ҪZ�,:��îv�m���K�ڿ���&��#�l�ә��q�>D�. ķ" ��$�D���	|�O7����x��\Gm����H��Uo�\P�\}Y5�3�I��0[�(-��Xo����p�n�zw�#d�A��:VP�I/�a$��yǠl��ɲ^�9�b�FH3��2�r��&[�s�g+�����[�y*��0Dǭ�1���g�ܤ���/��lY�*@�����6+�-�o	�'3���y���)�
T��A�t�f �G2�3�(�����?����֌[� ���D��;G��|a@�uđ�T�́nj9�pr �C�Wox���_�r���hӓf�|=�L�C����d҆���l�9�W�Ǳ3$ߙ�<��L �u���qmP7c,��'���B�De#�h�3�Q�V߱��7�"X��ox_S��X����<�|�5�8Ev��X�h��}"�I<�D|Dߓ��K�?�`GU!W���<�;H��r���۶���m�����q��`2$��-	����%��5M��<�C�Mx��?�s����R�C���0Ք\�,TGNXUk�%��#�ȯ1�t	�(�|h��X��B-�����(/��볗�x�	l�ASZ_��H/c�K����
%>��9
�*�͖��:��[�����aG�
���A��uV�6��+R�����8�A�̢���#|����G��]h�!�uP��iXy!��vg=�y*�TY�#B�U&I���u8�ul8�[��#�1|il�Ͱ��o/�S"����m���	O�MBb�Xo����)C�1�����چz^gIn�C��c��#�pG��I�
��N�kx�?�PYE�q���C�X:���q��P��#�p�,Y��-� ��1��sp�iL^����]�U����L����̯��3Hz?T�����k(N���bT��|�w�F`j�ox���,���|���b� d�F�;9[m4��
���h�" �,"}Q�"=J��mm���^T[�zF ����^_XgJ2I{] k<ڨ<a	� ���W��KI+b���)��}��T�O��U��o�4QE��ށ-ʯ��� Ut罹A���t���=j�=рv�կ�5,Cѵ�?��5=.�͋E�u@�V��8=M}��^����-�V��l/���L1�� DZbV{�A�?MK���g/��D
\1�x��cg�
@�̠���Ʈۑ�މ<CM��;���o����
��O��	Ї�#Eeob�=�s�%I��a�o�	^���{<����	jI�p��=D�P�+���E9C��σ�����B7ݨGqz1'�ӆ1��e7��/E��Pu����/
������0��}1�J����N?�4S�=���>!�R���xU������� �Y
�C�8.Z�+$�;%h��Y�N��`����
|�L��xEznǎ`y����E�V�J*�4O���U?��h�"����cWFX��D�ڼ�V�\���H�|�v��䅅<(:K�v�w9��-��������<B�B�g#��:��5ѻ�ׅ���=r!0���k@o�F2�
�$-=�P"WY(�@��)1{�b�Tx|օ|ţ6nM����J���V� �?��8�~�9f
CG?���l~ѭ煵��8t�EL�zxЖz��M��	u��a���Ą�*e��J���L�w~n���4�2����4#�.����7f$�c�l��hb�|���r/��ЗZ�??��M�l��E{VvRj�R�'�,jY+�ࢺ��>u�lf@!osC}��ud����4�ޓ��ؿ&�[cY<�����ʿ���;�۞:���Ps~7v�#�L�i髂,o:�K��U�9����p���(��g`1DP�%��#�-�:��Ө� �J�K@�k�Z� �;(�1����6����0�{J�X.׉����P�e�-ِ�~ҿ ʂRKJ��*��،������nr���G�#/���=�f]G.L�q|�*��	�<��,��Ty���Rf���̬u)l��~hT0�o��).$�8�� �g�q5M�k�JF?�%�-Pw��0�rBP$G��$���Z/�56�Y�n�O���(����WA\uЌ�]��WOJ?{��#�v`%h5o�mݐ��h3��@'���7_@��c��.8Okq�]��j�v�^I"z1��QΘ;�n��KǞw5ޕ�T�BE4�_���]~
I���q�>HF�1K���z$�J*1��$�}����H]�S�Ϙ:�B:+����p��us}QH:ZY�K�G��`� �����dZ��T�>�G�t�4u�s��1aA��r���OMW�~$��5Mii�N�����-�}�����3�B��m���f9��@����}��eln��0�o��@=ϧ��Pm�V����I��W�p��A�)�����Ѐ�b���Y��<�mڦ�T�%hr���S�e�e^�?�$ϩ�K������&B|�H���T����'q�� /�`��(���Y./�Xᔉ�qh���g;�4�M���C�����'^"37Lܘo0�@�!����ٵ7�R�FO����>�[k��Ҧ��x���A��X^�R��YD��?k�����	�߻�6��q��;!����v�)����c:��ƈ�͜��+�?��FX���d�;}R|>��dU��f�X���%�u��O��9����O�B���1
:��R�؄�s8����/�m�44�P���q@���v�m)�_u�v���eT0A�M���H>���$���$�xtF7%v4`�{���`)�YNq��2ub!3���:j�����k����gp[�\���x�s�0���������ҙPoқ��
ILs37O&�(z�	�љ��q�l���Vұg�,���w�����J��s ��̜�y�yrm��L��X�'-'��h'���l�֠����j�g���#�@n��x9�<x�������	{Dm��WR`�\�����<����KW"͎fDiщW�yG�'�8�|��ʲ68�<N�{q��Ӎd^��\���-h�K1�L���Q��8��":L�ʕfT)�����+S�VB�
?uiG]����ro˪� �B��A;��������l��n�O.42�k��E�#%]�ѴxEYb��՝yz��Qj5�v�1>�2��׼hM�7��9�&r2k��F*�o1����{z�`�*ph�z��[�PT/��M��t�,X��V+�iz��/	w��T�*�`J<@�A�v�SMSm�=7��|A2 Q���������ҹ���z0��>VP��S�1��|
�s%  �u$�)�5��NS��`=��{�ش�J?��J�����8�W�'R����ҒO��ș�v�|�7��>�G�SK	P�؟��ڶ%�0Kt��I��� {�2k)m��q��
�G��U����Kzw�!c^>��h�d�d)n�YuL� ��:����iL8=��0������Re��׸w����0I�(4���R��)�C�)E�>+��,�P�����F��ԑ��h�B$FJl����uh�K��o,G������n��a��W�� ��;K�J�L���L�v��Nn|����5e���쑪 &����{>������B_P�c4��ݣ��k����yЁ�	=����}�L��%�ɛ^�C��z�����4�����HX}ј�X��밿�('�߄���)w���Ҧ�1�`˦)j��^�]��U�a�����M�G�AtuQ�>lB���p�}����9�Ao��]�������g$���QY\d����H�0�DV��v�8͇�]�`�i�/�x�%u�Gw�������,h(�]��|�����0���
�>�������i|�!2	��T���r(�b�y5
�;��b�W������xݜ���ԃ7�OQ$x���I\�MF�
I�g0�F��+e�*XJ����*�|��y�uh�Ur����] ]ڥ7�P�\O��]� �F�)�+7͎5�&�?Z.�YW� ^d81Ҟ�c�[�	
��!���L0Ħ\A�h���?��AI�v��K�ˈ>N�f4E� bU�
�>P�.4�p�~|.�V.�W�j`�\e_�0V�8fd~�1	����G��h�2}F�B�_��1 M/�6�_�/0Ծi�L��x����KO4�&�'B���.kc�;l�]lHkف�7N^���m/��?m���l��;-�ߔ~}��NPv�qa)Xx�jA�B��� @��!
#�lk��i�p�24ލ���� �-��M�R���:��r�Tω2�]&�.��P���vt�e�*��ެ�t�[<0�M�B���� Q%�r%��r�B6N} �� �Ά����9ٳ���Jj���r��c:,���"8��fU���:���j�Df����`RX��-�w��6���Ҁ�rT��<Ҹ�J�.�[�WX�IJj�6�fϨzv��*��� -�f޳�¨<ZZd��{�-=���2��,�R.�zj�2wР@�tH|�MǓ�|OE��L*�������S� /Zr1pcn���GM���r�׺va���ۙLr���%��n���&�ac�;�)t��"�UI��X@9�Z��Aa�U$�&�U�?B{\������g�A%�6��}�#g�:�*�j��$<�s�-n�$��B�#v��o����#��5�0������'C��N��0�� 㛡)Z��_����(
jA
I�A����
T����w�ZK
x��?�����1^���;F�LN��G�r���J߆�0���s2��D�oa�	��K2���k�d�C&Vقfv��S��8& �f�M���j+ttH�2����O�+?0��a<�U\T�.b�44�g���X��l�suٝ��J�-G�%�Q:��Z3��6"g���6��^:�ٹ��I����I2��W;�4>�ּՉ���R,5"@����޵�-�b�T���\t��*�dB?��[�,�/}�'9G�U��9���kJ�_��=�O|�\2$��T����}��Yhp���.; �p�Ʋ|nU�k�o`"�k2B��<��iȯ��c�CVW.�G����)J�/��l.�jr3���଱c���gH�8H��ˣ	�H]Ԩ~��$|!��To��ۚ�����5���Z\��4�0l(vr�����u��0�"v�F��a6l�ʐ���a�`��1ёG��.p�#/%Pc���r?�cW�v�0`�R�iU�`(N�9K8�1�:��{�*���πʣG�P�dwSd.��7�ճ����Zn��W����}��)-k)Y�v��ؗS�a�D6�6\lNW���&�Ȥ�ڴ3-��2C�u���S͏�3cU5�)v��!*p��S�o۵kBf^�2�WSris��$ ���u��D}ڡ��z>�@�E������=�36I��Qcϋ|����i}e���|^r�� l��j@��iXuo�{ ?�h-rQ�(�(��V�u|:B�c����
�R������Q�e(I!��֞`�9�q�t(29Ze(
�/#��6%��R�%���6&�6�q�I7Z=�����$wh��c�(��Φ��4�D(յ�׍^A�wū�v�x$qI�蟅�0a@�(s�#����P/|a����b_�F�b�o����.�M��2�{�뻾�ʞ�[�zp �z&b;t<�����4�9�6�c����;uzXH�	\|F;�C�+�3;|S�[���fH�W
M0�Vߺ�פ��@�������:�ӈb8*q�7��mf�
.]ၷ6�=��U{�!�A�F���^�%�XU�yL����
j
�OV0�n�\>@6铃BI��+���ו������ @�[���6dГB�Q,߽>tg��Q��;�ry�E7�e���S�2�I����p/���G�1��^C9
��TO#[�_ǂ�E�\G��i~;����Q/�
RZ��[���*\0$B�>�i&;�lϣ���4�_3�WL���<�=d,f�u���r�d�N���� _�EKI����ѝ�����O����Ō��<�-H��E
���P�_��L� � (�6��{��� ٰq���ېy���4���w�y�q�����Ն��:��zņN�z7�̞4�r:�Y
�O�e���bbߞ<�j4���F�=�y"���^�b�(��E��3*e�tem��xE<^�:��r����]H���h_X������ڭ�["�F%h��t���� ��2���Կ�v9���f��ѻB���
��K8�%/��#��HM�3�d��z��S��s1E�6�eH�M�Y�N>cf��ci��=������X�_�Հ�{ߞ	�Z�[�[j�5�32�m����w���C�R��b��|��ډ��5���^��6�B+N��3刣l9�<����Ol�<.�a�ߟ�aGW/������fU�W�v�~H�Q�=吏=o��Q'9�|n�-^F����l��;Y��������v/v��d�e!�Z~���ӨFi�*��E�v���K0g�t�z~�J�d)7Я5/^�}VO�9���
�'=v$%�#�wy����Q��7�`����$`��u�%޶��mT�{b-�s�v�o��d�noc�
l>��d�O��7�PE�W����H�gw��p� K:t�?����P�N��}�#HeB.���Hx�0�_s��3Εθ��튊f���H�����tR�cs7^Hf�� ��Ƚa	�1�"/N��X��wvܪ��b�Qk�Į}�]�uю����e���/ԙ2@��i6�s2<��D���mR�7_ ���8Cv��^�4����^���8����p1�ԫF�ӝ�ݬ��
o��Y���	�4k��N��S�k{)��$e�^.?w|�@��EL���!;�?���ٓ(� ������b�t��Y�:���P4\|�Iƞ�*s��>��;.r���m�3hY�����6� �Z�E�#!��G ����e�2c�呗����|���E$o����ʊ�
�eNv�//�42bw	E)����F��}�\zv�a@\�	��o��%�|sz[�RVs�˰d�0l��`�Y�s���Se�}�=W����WV6pE��Ww�d¥�gF��dd����3'su������/�K��anO�V�!�]氀��_�󈞺guo=p������B'��0�B�?�QL����q6�����9ӟX>g�����
Q�e�_�qxϏj�\F"���.�\����J���X_�iMbsޘ���%�ͧĘ�Az�%��tÈP�މ���n���B�x ,�m�2���B�_��mڣz�����g��|VPGVG.&���� �KQ������(lF�h|����x�go:X�/JӼ�Hya�[<PGed��w2�6`�H�!Y����"ۆ��k��J3^S�}�.��;}��(/1����#`���ciDj�:][fb��7�i4v]�ƞj�����a��v�Ԙx��=�C9�ה���[����_���5#v�mx�X�#�B�l2���g,�};���$�c�R0�ր˟5��p�����D,"j_����<O�����G�oq=g�G��1�t�4h����J�>�wȐß���N.ֹo(��B�f�@�d�ہs����6UP&9��J�^��*�"'�V>����]���Ճ�]ҕ2� jM)�>�V�&�~ҹ�C9�՘~Ik�ǧxC���ϓ�%OD�����@���4���<͜nEm�����9��m�L�g��o�f�Gg�U��h��H�pu�۾>�&C_�T���]�Η�O�em��9������{1X=�G�D_��5�vt݅�ga�`�G$��;����5D��KC����coU�O�iW��-!�y��	`�DE�|�q�NS{�ƴ%�����<�C�BG�dl��&�� �Q��;�����7�P9��7@�t���p���D�
̆�1'RJ=A||D%	
V�\L��[��f��h��&Yp �Vi
f�W�U����N]O�/�p�K�kj���D��%����x%)�r�8?p�{�G�T���Y�ɶ�}u߫�|o�s?lL����,ߑ_Fo�^��;�=\��r�<��h#������D�>�<n,K���Ѫ.�M �����ڂ�d��oS�\��`�a��F#���tg�+�bC0q-1��[�-���:� ��Im? w��o�P����p�����	��~f,d>{ [`̍w��B��h�ăQ�MC/s�2�1K=��'R���H+�!�eS�j��;����9�	�.�������bN2D<jk�u��Q�����"6�{R�p9�atG��
�6�[c#l����� � �?����!�}8��| �Ԍ��F����S�ML��;�+P����O���|LYm��䟠��no��L��=�1R�e�S�%��	� �*,k�	}���~�e���0���X����Mm�{�D�-��gq�9���cmS]3��R��9�b��Ծ/vӵ�[�dy�O<��)<=6!5���råئ�S�!Q1^�����q�H�*?������l��e�����m�w�D��ZQ�vZ�$#�8 ��hE���n�9;�:!�y!��ϫ2C�M�d܉���<���:�W�נix�R��湜5U������C\��Ť)�ļ�����@�Ge%��ͭ!吆��q�.]<J�rn{Y��"I�XcF�9�[G�j��|���bf+e����_����۟	��+���nu�&���t7f9�" ��q~����02hȂ$=�$�rY�a~�w�)����U�~��qUP�㍦>Y��2@{���_ʲ���<���V�:v�3H�l�wp�7k�r�C�Ǜg��IP%�W7Y�cӀ�GMd:��OA�뤌�\�z��o�08��[��7��ffs۹4��g{���T
=�]	�0�~��Ҹ���l��ܸ�>U��>yw<���r���E�7�){�5�u��:��Z\�~Zr�	`H٪�0�I. ���,�SnF�zL:K<l����[%B�&rR���Z�Jd��JaCԜL�����
�vB���O��ZL����P6�3-#&��7��+7�F������J�#P�ON���K�wj����y=�Щ	�l���م��p�Ww�������4V0(�=�h�.\�C I4̌a���&�Ya�0J��F:�X��S��"<جgkL�]�SgR���D���-�&���y���b����Ԕ��N���]'���wc�~�9��]��'�A�zo���U���_#͏K{#��a��j���
PyIS"	��Q��>E>�9aj�����E���Z����^?P��9��liG�Ix"����b��άQ#)�tiHK ���ᓎ���O�w�,�|c��
G?=��Wz�;�*�S,��I�Y�ؑ��)y�H�q���9��p��������Ɯگlcģ���)i�	��QYD�q���m'��8���w�6�>-��ݷ-�3g	'�4���(u���O`CL񺸵��f�i�P��O�`Qy+��uјӗ1�rq�W�	������ ����10Sz���9�Nm��{0Nk�zu�0%��^=Y$�A��� 6�ׁׅh�7���[��%�IJZ곢�:��-�x�i#ʲ����b�������91ڈ�7N�'��2��ϋ�xc5�6F�f���.�-�Ǉc��0\ PB�D��OɅ�۽��+(�1F�XW�ޖ$-��	�۶���#Om0�)�k�S)���2��.�.H,3�̅��ѹ<C*=�O�z�X�O��|7��$�s*����D�*�*����Z���i��YP�t\�L
'�E���1?XaR:��^0]��?�?G�^x��6��_�Ķ���՜����B�^�G��_���s�j[�VT6�l�A�N���h㥳c�n�mC���.�L�&~�J��{H��f��9���2o�2�e8��PE����ޙ�ei��b�P�G���8�l�U��3Kp���)��!{�P�9�E��`j1������F��n������ބ~������_7w\(�7��"UPo�|�|(q9s� H���UJx�5��x��U��ց]IPK#��sU�X27�#q��q�.�G�����ޕqgk��?��4G+Ͷ4]�:괶�뒯���/�,���Ði�d�dK��_�nk
���>���G�l��y��W��t�\W^�K��k�?��[����f���R�I՞�X4l1��UX'�����K�Y���5
���"����vȎ�{Q�@��ĝ�K����}o�W2i�t�M�h>��Nj���>��e��b��3�7X潝�(���ѼJ�f�G����s�њ��?���ڡ5\pM����l��$&$|�O���Rp�XlF���+	�p��T0H�h���"�d���|x���0j�0{s��lg��ǚ8C��C��񿀥����-�5u�8�0����	���o`�ps�j|��N0�����f��o�\��ͳ��w�X�!�E�@�a�u��%����t��+��Y-�B4�V����?xDO�������@8�n5C��~1�'�=�An}+��ϥOhiSPc{���@�&��;����8��ް�H἞ȓo��p���33[�_�|�B��h墿AҲ��v�+h>�זe�m�ɉ������oi/��hI�o�,վY�L"���3ԃ=s*�/���߯��AC���)�%.֥�]�w^�\�9JK���_R�|NLp�Ӭ���� ����)�I�a!NL�쁋M
�~sT{�z�E*CWߍ4x�8�E4qR��c"�s�G/����G��*���4ZzC��ZO�\�)Q��Ğ��~��6D������؍��wжN�V��V�G1OኯgM:�v�����A�)�����GƓ}f���+R���g@v���:�E�/!�_6V9O�7UK� �<�J��.��7s��&�H�ˢ�O�N�k��T
������#M��� �#����l�[���rJ��
E�Φ�ܞ��]��=��	rm\�	0���Dj(�4G��e>�;D8��QZi��/� �ƨ!���6�Tc��1{�6�C�y�aZ��S.�D�4�%9e.-a�M6�����H"���ք���ڴ{�����O�nL�����.���}�jy��y��	��S����55��t����� .K0q�RH�����g�J/��Wc-���iz:Fe����EYwB� r�%w7%�x}m�
y.�M���gcm�և��IM���,�ʈ(�$ܟ廴��_�_�XC��bK�7�ϋ/$$t��+yt�E�&��KW �R~T��!e�iZD;�B�~���Wt�:̓v�۰��)�a���tt
�!��I{�[�2�\f���:h#�=�l��=)�=���8[I�ݰ�%"0�t��~���4ޙ��Mb�&N���+�1���t������"��w�{콢VN{��z�e�۸��q�h�d�)o,��W9�8����(7�B�!���걋�����C�Z-uM�9�#p��U�͂��'(U��R��zL1��-�g�5V���X���!6�S��`������Bh�Xҟ<i�;|~��J��0y~�y�c^��7ԅ	�LU�"я�i"��� �%���s����ZaYа`j����f��0(%��V&FH}���%���=��M&&�%Y�T:e���h��F�6��lH�x����¿���4�[d�\�IݵL�<~<����V$\����[m���:�R�ѿ]y]~��}��,1�۵����EԶ6|��D�p-��!�(�(��^<��_iY������}$a���x�:�AfF�s<�4mu��^Bl�E��Ba���N�Q^����a,Ղ<FX��p����@�f	(���3U]�?��a_�ʃ�Tɔ��@n$��o2|���-���9>�=���|��zqtw��~���\��Z�S�+^�"-������V����O�3щ�9
��ἓ�ucd��1|6X5Pm|T�����t>�����.�@IN=��P��g?�M �� �t7��v`K�V.��-XG�T[J��#�đF~aJ�͑���ٚtc}:$�����Pल�Q��+�D\�ߩ���E�̫XJ�Z��=�\��
ns�5Xu�a�)�$�@n��#@�֓P$�On~��6�nnd�{��HL�b���{� T���3^��Z�#�(+j�}�4FZ�Q"3���zX^���y�3S�0�D���- q@_�f�M�w�v��]h��6��Q��q���j*]�<��#�g���km,ͻ+���>�� �K��{�����,^��i��i���Fq��������5�?c	�ǮT�[�p�QH]�i�n��?p�Ar�E�7�œ'T���!����!�ՂC��z#挠H,���k� a�C4�;j�KG�?�R�l���ҸN@�8������_;��} �'�)0I
\�a@�2=|���k�q07�+����5�b�<�tY��n�(��J$r!�äPm��Fر�7�S�ݣ^��-#�&O;P��e�ԇ��L��Ƽ'��]��0��jƀC���}z��<|o26���O��*��C3�H9���O���(p�"=&S>V�&-p�إ8N>�aۗ5�6�Ι�� ���mb��h��&#���:j`�S���L�8ŽZ\d"�}�)K��~�gH���Sھ����jesv@Nm���7lCP�ᾜ�;͢�bVoB�'Z�9�J��s� A��j�V�T5H�^�DTF(u�_z�k�Yg.�tUV���a�9na	0��\�P� ာ�o+��l�ԩl���z8���p��,:}W�"]$	��K
�_-ŚL�Fk��)��Τ�oIA�3��YEM��#�p^���p�LG��%K1���%�J�	J�-STc:�ff��������o��)P�e��0z��4�4��O��+�F�>�mC�!��-K�U'��[���q
�]I{����2Mb�O�%�lz��N�X�Z�־�-%���ũ�{��Z�\�)�.:]6��Sj燪̈�3s�\�a�{9.�+�Hu`��>��Ýsa��.]�)j��F_�#%�B�,����Ʈp��S�zR�]��������6�7ui)���+_�5�̘3[���v��#��n�S�Hi�42��������bfQ�m�f��yi���S�+��1�J��nGs��׮�UR���}O���� '��3�Kp�p�*�WA��Y�`"& �	���8�U����'J���ַ�m@i��5\g�&�C�c?��Uꈣ�V/��Vf��B\��u������\'N��G`Y a͏�����w��l=����<��Б��~��:����|8���*�$��/3'Z�p��ꀴi�M�q�����<OC�!l�^d� /���7�pJC��l�WYa=ǞV��V'���͓4gڽх�����0���l뢜�=��WR�-����TWE���gs�S���Tn��O�[�gO?{��mX,{{\��p"Q3yr��+T0Zv��D7a�RV��7�f��9c������=�C���sk}����TI����/Uǉ��x�5�6˰�8{Q�������%	��LV��}�dNH���$b�E��E����ΰ�+�Wh�#+[�y�5T>�^�"��g��2#D�o-S�u`fxA�.����P�jډM�������pW}(T�}��������i-ez4��]h�I�.�` t��}-u�F�*�^�9�A1�eµ֓�*` �J�\�h��N� B���t�v�ԭ�_�M�6����.z�ą�0AO}������d�^�'��#���G{P�\�i��Vf��!��
h�kCf"sç�p����Fk	S��x��i�:t7�!�p�Л#�&(�4��s�"� �����O��hGL)���ځ���� ���s`��"K�Fȿ��*��j4{�D�<#}��˕���WL����w�3�{�ꍣ[y"���3z"�)���Ә���]��ё����jqW�;�8)�<U���7^��Z�X�xvJ��E��]:x�v���.���i�"t�fåמ�R�	���Vߝv�܍�]� ֡!
��%����Yv4Y��ZH��ȡ8s*�����<	���5F�w�#��
2������ׁ��μ}�;��'f5��S���he���_�t��m�98�}�7�T�+6����Zxt�C�85�Y/�~7��-Rx��=i=0�j�p�'�1!�2KL��؍��ç�W�!�>�1�#»�PK�*�wᙈIӾPZϟa�)�j��Mp��=�
���WML��~�v���4���h���%G�yt����W�`�t�=/�8q��g�ό��2�7įI/-�u�pO��d�릏Amo��seؠ�	��r':��?��:�8H9�:�����Gk��[X�Ös���N���&�4O�!؂�(D?f��i]�n�20��"`��������.���_&��T�x����n�/�o�x�E���I��1�����N�A��_)�q	'�_��:��u��N�s������������?��..�k�\M�++_���<?��W���&�I5+��+?�w`�X���%���)0��_�<�z��9i����+�G��$ֵ@��������.4�,��;m����h������4c�;����x)��dU�qJY������RR��w�S:b���@[�+Ԑ��^����g���hW��_Pi�l}���!X�xx����8��XVgt�w����ӱ�%��i�^"�;qA6�>��f[*r/��Ċ�xǷ�DǮ�'����rQ[5�;�[��ܙ/y���$��� �5�@�I�C������ţ2vRW�T�?�$���S��=�\̴�Q��dP"d?f��k�jй�SN[���\�HRy���H��/�
?��HїWݱ�=9���S<�0U�4a�"'�=��?�����>Z�>�e�U�?���k�&	�
R@)�����.j桔	��mr���I�t��oʪ��;�d�U3��ՌwW*�>F��6��PƢʻV+�M�@ ����!�R$I�+���䛙c��ʥ�o-1tcFwn��3��]�f9�������Ɂh'�OU�W"i�n�'1+n9  ��ţ�>�j�7ټKŜ�w� e�)���oG2F���,N%���L.[�Y\%R^>�懥�8Z�p���@�-�8Q\4��N��a��i�};=p�����L��r�X_��=ay�u+�Q�Щ M��I�ePux��`C@�����>�9-�IY�7٩?R�P��M��Qf~'�`���:�,�j�M䖏l�9����p���t?O������'��F���Y�>Qu=��b7v|'��uL�����O�����o�Yȧ���@�O�F֏����Ffy�v��R���}QѺP��R���g-kc�����ޞ�/]zִ��J�4eʿ\`{	���#�"���qͨX]8�ղ�rd��;.E��'��٦w�I����%���T�vW_����:�@���^����\�yq%��X�� `�.��)�~ŝ���f��'JR 	�I����E?��X^V*�FyFf0�Z�8���WS��o'�-�µ��'7���E��;� F�\�0:���Xe��!�*}ͻ��9�l���>W�/p�R�0T(�^nd�*��}z���<����^�_MtX�/4���7�D�]f���2�[�}��߀�s�'6Q����ߡ�[���/+r�"B$ �)��?�MEl��5����[��M�wř�"�BP)��	�K#���G�&4�\ʫ��ܽ�	�vÎO��J"ρ�"ݩ!�!7�PV����J�c86�!�L��`j�Ǐ�yq��ܮ�����{������f)o>���ss���"�*-��؟���u��U{}����Aî��W����Tڭ��ɱ�S�,��&��M87�����5�R��_JH�z�oH�(�}n����5��fd�;�ԐY{��BĀV���{S�Qi�fB�:���~`l�s�K|8&��ZDx���j�8�)��u���@=,[|L�,�A"����L[�t��hqR�T�Q`^;���(�M�ԗ��2xB�$����Q>�tҌ���T�c�.�"!#=r�џ6���ՔMp�����F�Ec��TB�=�)d�c����Hjm��J�arX�Xܰ�'4��������q,=#�C�%����)����=�L)s��>�����ߩ�F����xsZ5.��Qm*�<xv�V��p7.e|�k��&�� ����S���p��Q�YZ��;{%%����Yc��&y��G?CF?VQH��;�(��������"�
#2�c�B���C���{�C��S�߁�:$~�1t�`u�����C��gK��S��>����i���/S]��'�Y�a���7��dB�(��5�aX����-�ɧ�����f�o�����y�r�c����j/>�!cY!����b?3Rr_���*��p�95\-L�����Ԣ4p��;����5�>MTLYis�u�tbT.��i3��U`����*��������8�V���0i�m J�h�/�N���9O���ܑ���-խ�:�.˷�j&�)w?:މ��O;[����pX+��f*��[�;d�cOŨFt�[G%2q���r���ٶ��vR��*���
���c��z���qmT5�s�m\�����W�U˟)?� NO��XH:Xe,�Bp�	�I'�uj+��Q�(J�R2�ua�mO��L�m��r�SfY5������/�����T�6Т��y>o[}�J?9vI�F�hf�i�fcQ�� �6�����U�R����
�C�d������ �$�zg7ꔵda��5��.���jFu�Rj%��y�C�=��= ����}QYxGU�	���x�l��.�D�sk��%[���F�=A�`��V�mz��)�}Z�5n(^��A[��
k/C�^�n�a�'��A��6�[�#Թ��ü��G�$����ihA�Q�^f�cngt�ſ�1�h1�~�.��:ڠ<��!&�H�|(_��ǢYjtY��"	Me�M���ȸ�^vn�ž��Y�kɌt����2�k}sw���o�j��b�}�U(�Nl�l�'�#�x��[�_��X���\��?�ތ�����9F�e���TƸ^݉ \����eHU� ���?O��@�)�ܽ]ń������ww[xH;�m1J����I�TEr��A_����(7���a7�[�j���Z9mb2ʘtJ.��-�S��ݟ��ki�����o���y�Ђ����}r�e(�6Y���Y������ǿ�4��U�f�Y�ss�y'��6�8���0��a��r�CT�8��Bw�.�ʳ�x_Pn.��-��_x̅�/�T�}��n|3�t�d�j�d�R�a=�Y�,�	���a����$�Ű�;uU�j�� cʥow�:��g�t��q�4l
d������=Y�G����o*���2Ne'���M��Ϣ������|g�?�T��k�%�F���Y�\�j�/ǀp$w��2���*�HmV������GȆ=!�#�5Z����y���
�ϩ��.4�5�=O������v9�HI�������&}��%]<�[���6��Z�>�ZB5 ��(�~i��ҜD��m�`�<RD��~�_FRR��.U��O�zg[�����x=h�����
j��W�%��y��&�������`HB�m���y��
EA7�֫@����x����d��-��Z�Km^f>�f�Ѝ{vXr��];�A�<�W��Z�|�h�|�4�䤙=������%�n���05{��ߖ��ѳt 326y|m�%*a���79:�&��b�I���'������e��t,�w�e�n���@q�-��J�eMH�U�m9�S�r^�C�<j�A��0w�X� ai>Vj
�Xr�_��G�1��������,��d}V<���^��d��+K�@�6LxT[���J�R���gQ�X����~?C��ӥ�B�d?��Z�"ﬦ�C��.���|����3�|��Cy�N�B|��C�m3�YQ�L�qli-T� W� �Rڻ7rsY�ϼKN���*�h��P7�)����X�ӽ�R�����EEَtΌ:����������	�Df�mhJ[�o���M*����G��Р����S���O�J����,�]�%�_��m���p-��"q�n8��0>��$�( ��6k9w�S�;9�� �w������0��ʂ��B�ݑ��5Mmȝ�����Wե���BI�)H��:T�}=X��ˇI��-�S��G�2��1�\��p(��4�L�ս"�l`_��` �GA�
Ku"�P(��&|���q���]V������ct��	a����N�4�A��K9����E~ǝEz�o��Jʶ���Z���ț�i_Q�\퍱3vo�r�8vP�C1�Hja,�Ȫ��wYo��]?�#�~Py�A��4�c�m��Ō.U@1�G����e<b���%�gS��%�)�n�f�wY�h���E�Ô�A���+��Ao�y���ܲ��y	#"���8Pq�b{&M(֟�5O�r�I����=G>�z��3�H���H_:��d���q�7�ό�e�^��B R����iw��Fj�8pG���|�v�>����L��+�ϯ�����gE������ݨO�W4[�tz3��D'R�3C!qOr:�e!�c➅!�H(���n��m]�m������\�ȩLB!�P���Wo�)����g���Lt�=�_�u�V�����ޚHpi�<@r�m�y�M-C3<R����n���yx_�xY&���p�\8���{��}K\%�ʇ��ܕ4��^&T�>����0�<�mT�'�#`O��ak�k:�����FU��N�;����g�qSq�>�{#�l���T���IIG�V��y���7!���$խ@Z6�V�,�O��ĝ��֡�6�n�t�_��V4=k��E�xT�Z�o^"{��oB��<;'��Y<j���"U��Y!v�X�c|�y$����L;�|UZd���<%�)b�,Sy
�����[����@p�c��=�3��pa4�8��i��3mb�F�z�a�ġ������#����� MTI�������	��9���Ӳuxc�k�~�(Q�.׌z$0p2���J�Ɣ�g�y�}�	�����7�X��dV���`\Ͷ�=���4� ���e����S�r3D>CU�l��6��=��GU �V�$V)MQ0V����qDN�E��&R��Lh?Vw�.���a4��ܔ��ZQ�ͣq�����"JA�/8����$3m��"?���`j
�-�)űȵ�����Ug�WƦ ɑ�X'���u��Z�f���;���ZP3$HH�j��H���ap�fE��	A�Öu�����
es5�f��߯r��S��$Y���|��`27A�t�_Y��J�3"z|�KXF��g'����jGS��-�!ݠcŝ����������?�jz�Sw���\��A�0�|>2FF��m��G̷�͐��MM�"��&WuZ0B���I9E�TXs����_ד��=�V�~�n�
�O�a�SEq<��U/5����<1��ۋg(��OF��p�
�Z�}MA��1�G�5�����DM~c�Nk/S���DE�9UsBh�Q����ZOo�ZҹI{>��V�\������W$�D�K�xs�»�-A��19�w�"^�RWwc1�ࠏ��k�c��w���r7��Jǣ(�WS�n}�A�\ϔ\��UD ��L/UW^Eډ'�VD���f(�B����(�A�zc��a��+��,B$����w"Eټ��\}�bEU�H�\c�X��s���ˉ7��߁�{L��'�b}�J��kM�����|G7a�uk����'"�#�VFva߉�>��=��d��	�9߂���A�v�k�\p�ܫ
b���)�*�!�i\ba�es� ���(���N<���o�2��������0�����bQ���t�E:��ճ���@sP��R��B(�F�9h-$ԥv�>�o$�?����9W��Z�+D��mf�����6�⋑�dp�U��\�̑�N�}�����=���hh�g`	Fl.s@G��c!�^���;19��-(C�Hr%M\g���7�t��̈�m�0:5���o�e2���'���5H����P�gڗg�SZ�Ik6���!��K����UE���1T�!���?�OAV�D�[���S�{�VX �~�Ԗ���<;c�96Ӗ����I�b?���8O1�
���	rS�\��	bY����Mk$����\1����b����`ҢY���n��V=cG��w��Ȭ&��&�r�w��o+Mɥ�I��V�x���Wg�4��ͽ�٢?zV饂cB
��d�p:���"̹eX��/��|�~��
��г_�gC���kA��:�Vk�BGZt�p�������[fSE^}ZIB���Q� �' ��3~�E�;�z�y9�%�cN�V��p� �-I������
�ʗij��"�/y^���/�f&��%7��tf�A3g1�52 M|R�ЇTA*n�R��������F���>���q�x�w���5{�;���v�)��{�̮��Z�kN�+1F1���RMg���+��J��ew"na��Yo,(��˗G�����0l �O�$��Bf����F��pT� AVܪ���oyڲ����F�m7W�����G�������1-������J�uy�Ҕ^)^K�I p�g����G��E�7*)�fc�R�}-R*�_� ����F�&����S������ߚ�q1���&�IGh��E�bт��Y�AMD��>��5�I��=��������3?
>G����'�_�� �:Z��Z;�~��_a(��oS�X.@sP��v�H��-�-�N���x�Hޘ�����~Y�~��n�Exn>�o��Z��Ճ+�*y�>1,4�n_#Z�^}��|xw��xp�^��=�ps�,@>ݔ�of�I�4h4[�I��T4&ꚑV���O���^�?����G]�Xqx@�B2D��yF�P�2�i �+��R"�۰��3ώ�јl?�c���^f�����#o��@���>���k\~�,�K�J��\'��e�Fe[#���(U����Y�-6l)
$g���5~�)�"MC�Yʼ�I��$k�\7";�%�Jwv�=@�V⺷����3n']mؿ<���i���Vn��w����Kw���)��I�֒|o��������}i��Hz��	~DE��\����z�'u�@B�k�KsV��qLf}�[4֞���n��xۉ!�s@g������v)ϝ�����]�?����q���Ջ������ٵ�RF��X�.�H�q9:��m��(�S���hF��\�aK�Lޣ�~}@�%����� �&p�a��?��ɆH��j���fY��4%��
[ڪ����g(��d�H���\���ӳ:]��xKj-��8/�3����aq�r�y=��U�V	�p`?�4�0:��ӥ߮1&�7TWhx ��ji=t[#�pPZYG	����R����l�i�]%�	u��?���%'H��ߊj�6TDT�˛�93�3z��N�CY��I�����'AψVzVu�W���K��.��YCf�x��S<8ɓ��)2���"�_+}��{��C'�1*oU�ˁ^���^2�R����fn�o=T
�X�Vυ�P�}�l�@�=���R�F7�H��mog�17��p�{��w�m(�^I���P$Г��K��d$�)�\�gI1���0��pz�x�3w.O�A�yo>�i>;�\w9�!m@/�8m_�N�ܑ�"�Q�{�F4��Ie���_�3����������#�`�Ao���. ����j{]9����#*8�P��{�Q����+��Y�|t������Z:]u@��Ȏ���X�gN��	��^e�W�����P��xb0�*&w�Em\r�V��ez�V�r7��g���(�1��X�AG��1x���)�#j����u��6b���r�Ǆ���m@�2eH�{\-L����=�1"��vm���!�j8Od��ە�[��ҽ�����YKE �DO��wp�K�0��`R�4
ғ���KV� \�M�W�X;�%���l�v�9(���5x�ꖆWex��5�6��b �e5	{M�\�������FZ��:��Z�]�ϛG���a��;S��ر���J����ʻ��N�C����`p��-�+�l�v�Oԣ�?!KL@�϶Fk�#6�6�.�nU50.V�-{'f�8��a^�����=dr��jd��~�k�,C-��SIdv瑱�s^��}MWCϠ���bG�-�z���;#~�~��>$��-	�\��2j�)�I�r�uw���P�$mv������e�U��ɂ���П���Rv=6�7�Z�̻�Z'iQ7I`���J�_J���l��|mZ�L+�?����%�_e�7�zrI1��\'�+B�[5��ϰ�7�'�vKPS�P�kͿ�*R>j��יä#jc�(Đ���]�q�VC���G��*� ��Z�q�a�(�u��ҹ�D�s:`��r�2Ӵ�:kTb
dt��0{lD՘�/db�O.�7Q~��k\�w7�ҠU����������5�C�GJ$bD�hR�4X��ؐ�fǵ���x )�#������Bi���$Eo��\�N�M"�M��Vy�;�0�q�Q[+]�/�heK+^h�������.F7g���`v�Q-Ŵ�l:y�-!-��(�d�8 ��!���˪��������W���S]{ՠ&1��$��1��`�#/���g�~�T�s^cX����uM3ܠ�c+7=�|���	��>qHS_�4��G�F�K;6QR�Ӻ`'�k8gkl[��q	�e�����k�(�)��3���]��$�B�Ѕ�`�3��p�K�F!i�q�jU�Ӱm�̄"��얏�_�M��EǘD�9�MvS�oSy'%�"��ջ�3Jp�AXR��������\�BU@
;N�������n^��:L��������ʕޚsˎ��`*Hr��m��q�_�Gx�U��	�s���/K���h���g����Iێ� mQ�R��~�B���XXiV�z��6��3!ff�Nf�at�l=��Um-��v���k�a.=w���B��-��R_���?�X��������n��O�*���L �l1�^s ޽}�{��#��M�����l�G��H�pU���d�%���Rͨ2ӌ����Sm>��a����klc��a� vM���؂_~ =�5b�٠%�4o����
��(lߧ2䓧���-�m����
mwXN2�9�����S�Ga\�����q<�q��E�;�$��������S�h���mrW�gǐVc�?�O�B�(T�H������fd����}���`�l�6�=H��/�ާ%�Xg�Q��*�H�f߈�f��a��Ū�ĥ<�2n�%�7��?䙑cJ��t���ٖ���������S�ދn�&�Q;�ȑr�L�h��g[9)�T�ϸ3t�k�Pg�U.��or��P�sT��)M=���<���ʢ�\�>�)Y����|����	-���Œ���k3_��"�b��nU<u2�2_���pPI*��E��d��Z��|�I[�;����wִ�$�g; �?�L$M$C����!z5+�#%kB ��\�K:�|�	VK���2�a��(P��#�G�8�cy���˧K(��HtN��^�����P|��oN�2��.��%r(�<�#{�n�L(�@�2��- �e)�}z������c!/}�3��~����I1�;��:-�Ӽ�aE1z	=o���c7m��YǇ���Qi����A�M������]���r,����� ���
���U�Nx�`�M>t���#ƹ,L�O/�?
�[�g P2���OԂ�D�]����C�3�g��)���}��S�m�p��c�u_�`�M5"k$�5��v��ʶa�Ӯ���=½'πڶ�wxF:����4
��n�/0�FB�����DG�li�X��|{�A)_��I,�OQ*�gk|:Z��W�c%�4M����wrs���Ϟ����P- 7�y�>cqު��>���ւ�0��Q5(��\�O��r��)����=����3�������O��J�׾Ψ��H/=�,c-�WL�B>���"���Y� Mp���a�G��>��U�54W���s��0ʰl��~&�����}��`���C�o�K��Ŕ:P("�A�xY��z��.7�����$'�iH�,׫���/���\�p��v�yg�|�5�׺��Vg���������_"���t�N�����d��  qt��~jT��O�D#g�]�O�Sş8@V�r���_С��k�V��e!�v �k�;��(>�v�3�&Ǎ ���R�9�{i���S�\Q�\�&$���d��]n����*�l���]� ڑ��zA��_��x ��~1���{���LR%����k�t9_)�Ѻ�J|̮���e�}E����YS<�S��Y�Zyi�L��_!I`�x>�F4��w]v^tX1�N����(��+���CA4߱v ��}*{c�|rY��x�6V�.JɌ���Ÿ(�xy�']Pꎅ{?˺�ȐrB�+��4՘�/�!���/�(۫�E��՟Yи��/A��xB����v�Z3�[�'��0�Kk/��jj�S��߻G�HS�����a�(���~}H1��֧�/��a+ ���:��96g���a~��U��E�i�ꢊy�kS�)kAP�/�Ͼ�����?%�K;[2.2�c��������%P+�۟3�
��r��CZ�%`�YSIj}�]�ǃ��i��{!�H+?�n	-%U�'/�[\��dyFxl��=�?���Wؙ�
ۗ�� �*Tf�d�;���W&ݻ����K"�M�);���P� �@�r�3p\Oq���ΣKz���U06�3��u�Jk�K��xL8B�TKm�"��Z�2�TN}����8! ԕ�a��
�c��W���~�a:#I�i��GXi�B0$'Gp��8k����g�LrK��%���aK�[]q1]�մ��6,w��ӱfj��iLii�dv��2}���u��荨�A8���7|���%��Wb��i�q����U��@���_��C� ��vD�f۽�Ϡ2�`ǟj�7Q�-��h�?�}�Τ` �u��I�0�G�V��PY��KL���HZ���՟�U*`C�1�B���֋|!݈>K��Ӱ���~h��*{�q��k��*��H����l	�n�=<nV�fAv�n�V�y�FS��yC}��D�4�#f����H\1k���Kv!{���m��礞�)l�0�1������-W�`Á�	�̶�Xփ��R<.R��:�%'�x낀N��[�������+��ɵ���{��4]��z�1nxn$ ��\�9���.��?y��&Ӣb�x�F���,� �U�һ�l�C�L�'Erצ��#�G<[��yR̶��1������a�y�G�&�{���C˯�K�1���O����H(n)�B�7�O�����x/���3*��������P���ݔ��N�ò^���s*5�Y���6��ԯ��tѮJ[|�X��k,n9ہ����f�|���z<�9n�GJuKQZ���`������AӐ�&�@p����[�{��K�L��cf����8rKS���"XFa��z���c��\�Fɵ���.Q@��b��-W9T\��F�)�|�G6�w�KX	�/�+�[Hypp�M�P�'\��ZpJ�W�Y��DH�,>%�g[MVM���b,e{��s����z_X����a����-����K��0��fЕ61D�&j������%li��j���L�>�� yb�R D�G�p�IP���q�+�[�҂��M��6�ٖ�#UPf`��&t7�W7� �j�#Jֆ��Pc�S��}�h�v��)�}N ��o��[��/p�Eb��(�$��=z���a��������5+0��C��	��-	D���
nMlRK��"���Zk������V�Rm�X޺�1�6:�6����ӱh�5Fǂ� {n��}��G�.�����A�%(ķ��z�R�L�f���=���W^k�*
��@�+a2����N;�N�j�KSF}��f/ �{sI'�Gi�C �5Ɩ@��S����O|�$Rt�h5���t.S��o�.��S������!�9��}��̄�WK^�b�pF7��^��y�f}�w%�E����HT����	S��i�0μd�j�Qk��n�����]|j����O�%�����K�lZRH�N��K?3~~����j���B��pz؝�˲�g��[$�-0�wd4LCW���?�j�S(�3�S�^^7+L)Bt�ɧ��Ç�yk�@�wsl�k��!�)2�6�Q��\~����wD}G �n��1���מJ�������%��ok0CVw�>������IN���(.=�e/���A9��ۛ4�?�F���$'O,>7��+Lb�����-y1��sh�bOt�]^/n˨��'
���q]�*�Z>��q�؛��ߣ���{���un�|���k�eZ������N�VY:��^v�s��-{�1��^L�a���3�'J��G�[�f�V�U^��Ol��J�  4&j�8����������{i�c�����?K�О�A��m�X��g�-*� _�Mp{��Y�8�Y��H�4�tS����j�qc�R���I�a�q6 �;0���
f��L�9�<-��.K�q$�N�3qG`W�Is@�m s:5�79���6P^���J�����C���o�v�$�فN�InS3�kc��^e˯3�x����*�y:��;����"Cd�%��o�5�MRY%��)S4�s��2=<#��2⟡<{��s1�u �	.=x~&3v�SV%��ϰ/�Ꭾ��(���pW����S�}{"eh��]Y�0�l���U�%�*\� o�ޠ��5G�O�_��ª�
�!�<�Be���g����$ �:��9��Ok�+g�9�D�7H������$[K�z��W�Ji|[/�p��ڈ:U� Ϟ��?�Kh��Z��W#�C�@N2?<��nn!}���J�:Ǐl;-�i�����xk�� �;�|�i�!�m�,͒�Cpx�u[h�{���]�K�f�j�W=�i{�i�5�n[xF����yē&׼"d��%G(/_4�����^-Y��]]J���0��k.]Z��<t�]߇�f$G4uN�3��/jT����$�z22jJ��U6bM�o��mYw>�u�f���̴���Of7�vd�@r~Q���ѫm�cX`&b5�i5���ֱGk����]",c $8w�׵��i ���\�@-~!Vh8*~)F���������ʅ�£���Ԛ�%��C��6YŅ�1<��~�h�~ܑow��@ӗ\%k:�|�8gWF�H�v��d��u��[JMr��Q(�X��� �BG�n�h��� z00�j�TlU�^WO�iW�Dv/�4�}&�p5��Yp�-!JbN%!th�*�70�m�����8ˮhK�4�/n��hW����[:�aq�kz[/R������ �>�u��6d���P��e���=Ӈ�z�0m���'������2�.�M�th�\��c������da\��*�M�O�p�`�e�{�ߞ�ϱRi��Ӎ9�.?J0��iqa(��.rsF�|P���4ףR�����t'@z:��9y�ܟu��[�<�h,H3����e1Ϙ�P�2�~�ˆ��=,oؠ�1.P(5ij�;�[��}��Y<���_�ԂL�3 o`1㐇�(g�0���R"���g��ݦx�<�������~X4p�(�6��Q�V+�W]�Ls��}�JlYt�Q !!�Xy?!5]��.X�>�y���S�IC;��S�ι�@"9pPF������i8\���2�����Ĭ���������Xs?��Xsi�̘h�/�s�S��V�$���>u���RVG}u�N�:�����ҖG�����L��
��� �[�Y���Q�{=b�g��N�	 @�W�_�b6����QWt�%�"r: �=�E�-F�&<p��UC��	�K����c���-�eqӘ /ID��b��][P�2]�5�p"��Z<������P�?���u�Ig��)�F+:�]�q����2�+c̳� �E�f.�~&�		~~%ئ��n��ؘ�B؁�3�:]�D�"�'�}���l�Q���q1���=ˋ�����)/�ɏg	�NO�T*c!��$���@+�41�r��%�z)I��D&���;~d���l��D����Z"��Ԓ��H �l�pF������N�;dܼ��i�퍃5�z|����u��aV�\�������iqa>'|?9��L��dm�?Y�n7QfE�6E���=T��*Y���@#ӟU�{�������-O8��������xaٽѳ����v%i��dy�fBk�E�(��-�Co��8��(��7����0�M޵N�g����,e�7˃��h(�5	h�ے��d��|��D�u�Z;�R�r"&�WZ�֓vc�4O	Q�>��~Xqy��x�Q��Bi%Z½�^a[��{�PK���]��dQO�7�u<�PQ�V�x���t���L����z�J�U-��8��B�@��٘�S6�z����c���HN��l"�u�'��S��Lj�co�#Ku���T���K2��wW�yd=�NS&�*O�s6�>�#����ެ�Rn�`�|=���q��P�p=l>$����%Χ?��/u�h�3�c�Ibٻ,�ۭ�D�Y��{$�H5h�[n�nv��^#vA�e�ʟ�kj���F�å��r.��}�[�:.�B���Թ�'IV��Şm�;���J�����n1�R�	�t�_<��1�r�*�B�i��!�Dd�0�kYo�~�.0��N08�t���	΋��4�Z8 �W�	�y�C4!�P�|晉�z	��>�
��DdB`���8�ϋ��-�ts't|���k��k��� @��i�����w�*����`l�&��A��m��aĭ������>��탤����M/֠��s}�3�f�<m�k�İi�r�4��.�8��Ya}�V~e��9���S�^K(���['���hd
���2ulM5�.�ē6��I\x,����d4��Ah����Q���7*K$��ǩJ�K��G2���>��e��S0��ސ�xH�9h��ϕF�� ��R����6w)�/<������><2���K8��H�b����(���&S8�]y��/׋-5X�Gs$R�'=�w���͵+qU�����eUN�������rxԠ2�~HG���Ɗ�&.	|<�J�I������t-8��)l��ncRZ�ܪ����;�T�ϭH��B{:n�ى^�	c�x'��c�'JF�s���� #��{�鵉K̢0'�/ǰ�m{飏<�ë�QR������5����D X�^��g��j�	�8λ1#.t�!�A�"���&u��U��j ƞ,�����o=�9U5ª��2���68dgtB����`�����	�k@M7.i�������E6iO�*\9��~&���E�8e����m��$O��V7E|U��E�X9E���Гt���R��V�LA�s<1a#c~ͥW�6��3[N�ޥ�P���v����X	Re�a��e����*��l59�=�j����§r�M�1��x ��N铰J� ��SG�Op�3��5��We��G��T\?�D�&�{p\#��P�8������ u`�ci�]�O	܀�.��i3��Vοt:�Y~�;&�Y!�^_d�>�e�JcY��I���]5��</������Y�0���u:�+yDB84��{���}8B��N_v>�����i!4�t�P��[W�1��޷ԝ9 �N�lY}Ʀ���dJ�V.�wP�a3ϞF����Oe��L3r���9�Cب\ߵb�C�*G2i��0�d'E�i+���05�v��,�����o�$��x�_v��	�yΧ�KM�σ���Ey�
��μ`[�S��)���4�����S:2@䜔���!��g�"t�6s�>I��T�8:�_��^�K�!��ԀĠ�Ȑ6G�Dgń>���c������?g�ղD"=W��3j���v�ZF;��TS:\�v�h��Ű�d���gm�����]��������5:�X��[�sl �.�#���&yfw<�H�TD�2���n�
>Cd���R�M�<]�霦��7}
I?�!�������|�h��Q\%�]�A�8��zي1��o�1��W�nq��h~�Ћ��&�\OB}1��5����nV���P	/<��̞^�m�3��[�?l;͆��M��B�'5-E���pÛ�h*K�WMc��we]�P�6�O{��6%�]�M�T2C����tg�֟~.�*>5*�R��"�����y!��ڊ���>1�}�hR���ӕ`�$��L*��o�q�q��.D �~�: ��ӕ4L�pœ���3>ꆌ��|UE���X �*#q"J懆�(��i�˪�ϩ�Jll��UZM���}VI#~�W�N��\ד����������0״�V8��T��\�a�R����e�us:��٦n�������=�g[�A���>/p*�\
3�f�U����k2���zC��őB,��|6&���4\/�,���i��v�0��(�A-o�(�����'��"�C��\X��
XW�A��PWwL|F�z�������~l\vE?��lE(��7]���C��dĕ��7�=��j�Ņ�4����P��5~���ģI��ګ��󟑊��Դɴ�+{�#��ƨ�/ s�DB��?��i��D`�qv�����������u���2,vY��H�̱��#�� B4�g��k�2�����h;���Z�3~�|���E|Jg��|�v�Ԑ�ْ�j���H�^��~#�yJ���,�����N����9u��'ÖҖ�B
C�ڨ�y���. ێ�%%`�e���`�0�U>��k�1U�_V�|B칟�/��Ҳ�1�������
K�����W�����;�E]����K�t����7����Ҋ��������/0���ƍ&�0����"�w�+�a���#! 
8�L���O����Ǻ��`kW?���Z�����K卣�XvO������@�1j�`ݶt>�\y(r��[^r2�+΄/
���@V���P��L�YO���%��zE�Ɏd,ٝ>ZU����3p�����e��Z���г�p=��:�fs�ߛ_6@���MM��y��נƴ�%${t=��"LV��j�PӐ ��%c�ќft�!L������g'�1�JP�$�����k,���dE&����[���_�*�cyq�=�T޹��e-��SR��oS[ql������S�;2o<��B��E��b�TV��R�R&����,#��^C੘���2�M`�.��q;���=<�p��.����n���%��9�&�������[����m�=�p0��Tw�!��L( �.�Qu�g�3�^H�4��p�NJB��I��&�"�.!��K�ѯ����]A`�0����R��8tS)a��uBM��=HC��??��k��!A�R�o=s�jPcb٢œ}�Gz�(��ڹjH��Q�h�(���n��D�Q>��f?��#��^�&
FFvUs��t��im	|�#�_����S,&�n�֌Un��U/
�J	���Z�U,��ސ+*�3)��=g�Gr�h�[�yR�哝i�?�r5��2�4^n���˸F��n�z��W}zM�{�%�����J	A�݅e���7�J>@	W6����>�.d jI.7;�����D $���g*��FT�}js]
��6��mʑ�w���ֶggE
ɯƺј��FF�d�vQ]C{dp�R2G�sD�Vf�
�j}���D�,��@1�0X��_ODf�;��@}ǌӛ�.�G��V�}����4�Od�ĝ8�v��v`=P-t��+i�����/M�&-�@�'�0?p$DV�a��;2�y��qa���DeĻ�H��2�'J�;�oN��`�PJ��0� %�fL0
f�;�I!Z�A���Q5��o�?�Pr�N�21n��Z^�M���k��"2�-Ź_V�~����b���(�C�`3�%@<�r~��+�5����~n�'�ur�'�Ͱ�v9��p.���*r�K���.r�8�ڟO@ڡ?rd���M��^�T|��k��R�!��/�]�,Ӄi��ߕ�����d����ō��5�Lv�baG�����<�c��иzGu-t
�)�����Ka[y�e^� ���"����*��l���KtEr�5�F��a� #kS���<�A*���QV�]h�=�m2I���܄(�	�b�9�+z�O;��3/<.1��z�[E�O�1K�������Ht�qjr몄M��<0�?��"�cqn7�ج~������Ͷ;Ad��_λs���<V���
�E˱�eD�����c�F�pJlv�R�;�]-�z~��k�ݼg?J�85�c���5���� �V�󫎽u�6�4�v�w��V��|����fS���`+�T����o�H���9T��G���#�2�9x.��F���R������X�y23�=�C�qt-�mdWT��©�<��<Y��=q)C����'�!�~�Bm�}=��Eꠥ�揅��ub�P�#1WĒdaw��7���]I�gG{/��=+�i٪����ezx}M_\���Pf����u��<����s�t��S�ӎc��I�y2�7&�IGgPc��/�v8Yd��Z^��P���|�L��m*G��PE=�(��C��AF�o�"�fh6��ݴ��;ED�{ &謱��Qq �?��~}<O�T����O�1�Q�
!q1a�uqs�]X�l���d���O�}��~�zcF�
�
�	��j��Ϙ^w^��ك���v����:��mD���0��=g_N��M���58S��� ø�y�)�ĽN�Nj2\lVn���V�K��V���گ�@ox���c@�S�YTi�MÜƂ��Uw��tS,�<DL���Gb$d�u�åI�4�<!5C�� �>�:�"k�����Cp���!@Y�ψi�xXx4�J�2>Ҕ����&�x^�p-��Q3dF�7 �9��1��Nu��;���]�ْtK�$4]�D�ΩzΖ:*5��hљ�X�P�Xi��ٖF�j'v���J�h���J�_�M����"_�K5�9�Zu�(�U�#k��� ��j	���s�����8�F9z���<gWt7�k�F!���L6v��b"����+x}��|K��	��J8V}��qUJ��AOar�|l^� C�O�фv�sY> ��_2��3@#�rR�]\2)$,D�:[��n`����[�VeK�o~A9^��+��2o{wGlB��V:��u
S�M����CI�����Ķ��@+�}8�?���E�|ڷ�L���7���W@F<Uql���]mG��7d�=���>��z��Y���Z�:���&�q�2�2�٢�ś+�.�(e��� .��%s�4Ϩ(��<m;�I��k������C���Zr�x%�<�C.��Il����5��Գ�V��,o�x)y�f����UUO*轔���8�Sq�o�jN}��.��M�
���ޔ�y���3j���G]Q�������a��@��q�M��i�����a v�2�c��'+�fe���\t%��.��kN�(�=B�46����^�B����4��]�$�	��X%�ɘ=|�ae_䟗���L V���T���o��@�I�{���,������K8xSa��O��FHQ�-z��:0;An�>x�����N��'~ԓ�KKS��2H�~�0h��Ӷ�J�3��w�����V�+���.�΁��j���2P
�r��Y�:�N��� ���Y�?���)Si;Bh9��B]h
��cz�ܲ�EtG���E��XQ�0F�)��j���K��qЗ),h~���܌�d&eq,�9pt��z��wy�7�n����	��rU&= Ft ��x��=�.����:��L@�m�竌�����C���A(F��|�p\o�o=m&�CV���u����jn���t:O?���!���3w� �|4m��t�$?yZ؟\��K�i�oB��*8rX-���M��*d>��r?���V!�}6c��}�rr���[A�ޒv�@�
P���X��;�O1�7��lX���9k�.�!b������ E�wZ���I<$�[��*��C� /Ώ)v6ʨ�`9��Ѹ2�D�f��<YN������h��__�5F��/U%r���;l��6%;?�����(#�:_�џ}! ���l?�;7_�]�*����y���8��X�-�#��H��rS�Z��n�՜`'v�$��L����W��[ic�h޽g?���r7S���~�B
3A
6��0=��>�F@�V������Un	D�Z�~Wa��~��<mx��H�$p�d�s��p<.W�(�.��Ƥ:x���b�_q�)������"E(�? UocX	֑�>%Bو��<Gd��$���ʔB@�A3���Yg�^JnbZ�F2� ��{��`X���*8�DC�aC̜�Jvb���)����o�v:�[a~P�wKY�<uW*5/�i�}�S�������($��[y�r�U����@B�V��n��k\mu��짶N��Ye�߭�zz��a��rZ�0]&$vTM�|�b.8����j)������:��OZ�K�҈�`�`zõ^��E�h��=
�,������f���/�Q�ĳn�%N�}$���pW�8A���ǃq7�ئ��u�?�a�̵������d쉕0��E+>�t)��(S����y
�#�5�Rb"x? \µ�̈��'-B0'r�ba�����ޠ6u[[dS���;�Χʖ���Ĥ �H����t;n�'-̑`�u[� M�7���v3­���]6g�ŀ���Hg5up��hf�i5����d�����{�0e�C�e�� � 6є�	w<�mh-*�5Q�P�D��VP���"^�c�O�����̡7\���v��b�ym���e��p�lF��J���K#	�����`�L�W�����[j	��杶�,�@�qϿD�.o�qr�!F���L�E|� �ٽ�,__�������(t�)�H[�|+\�VT6�MaT{�8M�v��x��f��������d�?㰮���x>��L=G������K3*��d/P��������.�C�O�^�L�C%�]ϕ"4tcx��������i���̈���j��\�v��,Dγ�X��o'y�eK(��-L?xb��8�z����(�=k���ʶ�ɠ���>��+���SoL��uM�!�ڈP��+dIab�H�k�Sk�,�:,9xL"X'������#���&�.�V����-�(��lA��;'}��l��$5����Q(�a�1[â���B��:�CF�	dzD���n��Ŷ�;6D�W\9Z(3bmJ%Rb���ß�<	;�ִ5�|�]n�l��(d��*��ϰ�_���c��K�?M�9֯7}���T#�#�����|a$�8#c��][�d��%�h�zX����9K��f��Z�?������D7½�¿��x}#�{B���9���8��l-�n��^Vb�J��|$�iZ�	�wy ^ϫ��pӴ��V�E���i`��������]Ň&yuY����I��Uړ�^.QJ��0�tJ�,�ʤLozڔװWeE����4�GvK�N_�� ލ�'�L�Y� EF��ŨF����-5*Z� ��[��x0�>�gz�U�J�ت��!�gS�7��b��:.��2ZX0.z���-��i��}p��/��g�ZQ:��CZ��)��������<1e��Hj��x����=���Z?W�M��b':.,~�ž�j�����f����sA5��̧5S! wE��a+splO��@��q��7�����7�����߂�ܦ|�!��Ტ�m��+�:&��.�=ߴB��	lN{�}UE`�C7��t�Ũ�U.#{
�rB��%�̀&�g� w�Oz�X��F%�OJ���b�΋�mk�	k�wbYF?@��
��Pb�?��SV	eC{-�y�n���pxK��q��C��WA?'k�[c��-gr#�=��M��G%*���sʲo�e�4˽�=���a|�w���Po���VHms���miUxuf�c�-�g�*BC��&�H�uUO�5A {��L� ��䲀Tᝆ�>&q���\%�~7E��I�ƣ�\��h3�:Ex�f��K,Wr"� tLO���g��~�X���.�OϵA��,��T���k�e�t1�S��p��Ȭ�اh���"a�O��I� �5��B�<�$�	M���1���#;?�~a����������Q7CHu�<r��3�S����o�~N��>�~BԠ�-cj�I�4'� ']Y�C�*���Ab׬đ�E�bH��Mw�7�x��jq��=�K$\`� :-Ꭽ!dy v�r�eC:
`�c�.��9-�_wD�ތ����n�Aw���J� qޤ���Hs�n�+�粵oI�lU�8(��B?��k'�Ւ����w"kFR����ae�a�|s���>�j��R���soE�L.�,�-�?n��j�4��u�(�|a0؂>�>�6�������G�O5�*�	��c�,� �Ǒ��n�Ȑ0*v����y/�87�1%K��%/�V"Y$�'��!LP���z������mY��j��Ҝ����}����b�%/Qj~|�OL}H|���^����ǸK���v��q���<���K�:��G�q蚏�L�~$����]�㤽,?CE嚁ÑQ����n�Y۰v|�Gjs�cb�PLdc��!��
H�
</c��sz��n����ʫ*�{C�.x��ϛ��3oܭ-�Ύ����?�cFa� ���6������J*�z'"곱q͎���P$c��b~���:���+�io�l(��E&���'��n\A�9<z ۷��$��$��z�-9�J>`U�u��X�]Q����w$ ��&��!���}(���q��]pt_�P$NRh��5|#[u�s��X�A�9�@��!�}EI��4D��"��U�����'����˨lY�_�0����tVT��PV�nMP�st��6|Lh�E���#k��k���;�"�+X�,�q�V�J֚��z��.�����C�\������?�"��G�����a���<���(@�3���1�-��E-0�j}���"E�Ea��SJ��`����qE>�"3�Y�'Հ��!h5�I���;[����ޒ��0Η�І��Hs���a������$п����(�-�:od���μ�vj�i]|�����`��� *�D��,�He:��d��*h.Xѫ�O�=j~�v��cD���[8�B��Xo�����������0s*鲄����n|�k�_ώ�i�������aF?�$#4�8	�|�����_��_�����cm�����8e��;���|�9?P�^(���U�XY� ������G�ųrj�]���LIq��d� :"�K�:���X���l�!��܇��1�<&Y�ȨVdcXt���LU�=\�w��+GKD�����y�(:v���S�V��U�2��@K9 �KWJy�p��� [r6�'!n�ѴױAuM�jcW�yu����u�XYb����(5�|�;W|k��T�}Gn
�ߨY �sd ������L�؅�������01a��Ǧ�ew�����b�uHTIl��F��B�x�n���*?MĦ��JY����kf�����#��Y�}XZYR�#�c<W�y�p���TLH=Ѷ6���0Kfo�Q�;!����1�b�4��Ɨڢqd}z�Zf�;�h�pؼ��:��x+�y�<m瘿��x��v(�1��U��Ӕ#2�d�v�ݭ�	�pA\mQ���9k���O�K�C�HH�kSl�ņ��1����V��� g���7 ��w�ߛL��=g�I��r�p�k8f�4�����u�,��)��a��n��Q}����ef��G1i#nS��Q\�E��������	�v��(�2v͢Pq�n?'�)H�Zk�F����W� أ!n����0�y%�#�R�*�$/5C����<J�puW�QloVs�A=/��mzX�(F�{I(�Y+e�i<��A[֎&Zk���K��p��~T��#j��ԫ�b��f\Kx��>��� >+��I�S�����m��9��7*�I���RHq��ڊ��ԧ�a�6Ȳ�5	op�6��P�h����!y�dÞ:8��gv���f�cv�nMU�g�و	��м�oFN�V��F5&�z�M�;�-hb05E|ZK���^���"#�@�S�b6����|��	��UOYi<S)h`��>"��h���@7W{�1(ub>��C��7�+���&\�1�m��)����p☀�9��M×FZ�%�^���N�X�8�4A�Spu]eeIWn�9�c�mE���,�Y�K����U����,N��ձ	�y��go�Z���P������G����7'KB�`�dk�ݯ�n��{��gq�5p�@��h�v�� %�� ,�Q��q�KJ�%cG������W�E��g\L� �I��}�:��/�B�1Z�Ј;r��xfzMN+z�����Q9�����̿�B@��G�ҩe����Ⱥr���Bn�rmh�j�=w�Q\M���F��E�^2؎	y3�.˯s��}�ĸ��q1�
[44#��j��9W�����T�Kf�lJv��c��qqŷ�OṬ��낃����Tnd�U���e�Oa �tx����`.��a!�����o����^^� � zn���=q�I�물�{sj腞�	��}�u�Ĩ~7?`H��p����-^�	eP���a�Y�Z���1��fg���+s\�HHa��{O 	��J2�l`i9 �mqE��t�kg�����%�z��z,�\�)��[P��y���|����\�-�pq�Uf4�*�S;c�����ă����7��Ś���s������ �-�ȹV���[��X�$�3�YL�:�\����K*a����o���|6Sa��Nނ�_<�5G�6د���*����۞1YYeC��*f+Ʒ�j�^����B4`�8� �!�56^/`oLZLD���
|�-����*[�z��W����)���3� ��/eq+K#*^\��ۺe���@�<�HUR�xi�K�Q��$����HmA��y����S�Z�8cJ����/�_9�|嘜�\_ð�x���	��1�+�=C�f�q׵�G0ݢ,Q'��9f�?ģF�2�XtC	"�3
��*��G�FHc?��FJ�bӂ�#{��Z�z0��\���̰0�g�8�V�ї��iR\tu�6�����ii]����W}Pv�#x��8�r�)��|V�Ł�JL�D׀Ͳ!{Z�,���� :׵hTk�ə�C՛�7n�V����Ʈ2DjC�.G��a0Χj�7Ό%=;����yaZ���ԯr,$l�]��07�c���e�o)!�:��H��\���g��_����s���f5��E�o76��A�&?/�p��]�>Ik�H��?�d|����xDh�j���r��($�\���s�M���I�S}68˒�8ٖ�z ���AyykDBA�ra(^C��g	B�7�Ga*J;��6�¢��c�n7߉^"�V����ep2_o�Z+d��9���p�C��{�3�"x,5�i�#%�"v0�Ad����.��
�?>HL�#o���tq\0���f�z�b�z��5,�)�l���" ���:Fs>u�C�ƁZ��*��-X	p}�0bi�G
R���̛Ӫ�*�ܴ�9'J���f	����6�\��y&ͅ�!���QW{�Wl�t�贲�(+�W�V�3����4�����VҊ�#£�?W��F�պ��V�`XxX�!#P~��� &��Z q��E�]о�{��I��KKTT}=294尵&�(��ٿ�+O���ϰ���m$>�S��q�PH�H��K�-�ȋ�D��cG��Ƚ����D�,��@V�����y�\qV��[��;E[��r�&I͓_��u��B�ZZ ��o6�����3����5�=�YX\(���=[5(����.�K\��h���rJk⠺��K�����DQ\�s{��B�ڌ�>Ǉ_�}�ڂ�r��)����2��݉졕�w����	�<�2���<�og�]�"��ل]��>T��buǶ�R5��2��^��;��6c�Q��۪?�I�3.�^�Z܂��d�B���O6B����0}xE���]�dh��	�.Q\~����d���ֳ��]4���⤮<�S��ŕup�{����r�+��H��u�n���n
��Q��|4����>�=�QF]Q�;���l�� �H�ū�^D!���� ��T�s�J�65�7i< S�����y9�ӆ�)���� IP�3�~�j�|O:���&}����(�'���h-�nҽG/i�`��~�o:�F���������h�z�
,DCd[� �K�=���݉6�Zy���Jan�O�N�F�g�n���v�������5T�2� &y��.�˲a8J�'b��%�]��⩨ �J$���f[��U~9-�����[I�,q�?L�u�3���q5����d�6%�9��p�8q�W=�6O�Y'^�����e�ĺ@�+�rw��b��J�8�Q�?���~�[=�P��Ћ[W��
��~���ސ�7��洕U/ $	��"nb�~9�p���SY���o�^/&�H�+)�y�)��`�^sku��fAp�w{gpVk���t.Ѭ��A\���s3*:�+^2��&�o߲
�\5Sme��˫�Iٷ�P�ɞ&/�l��{?xrk$tU\Z�l0y�w/J�,�~<͆�$�O��3����/]vM���`nu�oI%���qX��u�L��X���rr�y,��2栩~�-���C6�R��Q�iڹ
�2��=ЃR � ��41+=�pU�H���������k*�O��J��ށ��e��!�VG�&�)���GQ3M�'UsD2��B�GN^T)`c���VS]�kȰc�#
�(��in��e�N��c)@�3�)�.}[���	��`�p ��)�'�������c���m��,�]��'j�s�ă�^}g������_Z�ե��%{Z�������N�T�]hGE� ]b���"��^y�Ɨ+��oQ�se�3S�p-M%i���`��H#@
./2�_��~���&3q��+���WdOT29Y��e�ԉ��*<C�����E�Ul:W��/�����Y�����T�2��O���y����u�U���"�x�����<V�ž�7L��w��+�考����s��(���_�/��;_��=ސlTm(�%$�Ӊc��vh�d�����]%�Y���g�E}�QO��a.��w��ZTV�-��p�����ؚM�9��/�|��)�O�`��pt[�Z����W����.�#�\���gM�-���qY~~��A�ž��i���u�=1j"�YM�@x��=���*�&\p�U@^g&���́�b-�pO��I�DMcu�����F�.�*tk��bkD��c���JEyP��g�!�H���GCL�����K�k?Z���W���PT�"Ǟ&�&-*�r�]�u��I5��\�"���}ܚ]b�<c9z& ��7�Wc�b�_��p�����V��]
��� e��P���x��=r�}�}4���
�M��������f��/��غ��͎cV=1=�h)�W-�:UZā"�o4ĩ?�'4\F;��a�^3��Ci��F�6U�����:7��1q<�N�x�.u���u�jFGi�拞��FX�-���o�>'
~����!�)ͽ���&��k���iW֝ʆ^z��v�XЩqȸ�~DX�A����~��\����ah�����������Y/�`u��߰���#~�B޺�G���r�}j��`���FE�$�,�v��ϣܹ&Y2��v�	� �;0I܃���Ǘ'U�w�8:��Q�D@�0���8ʻ|����G�݈p|5^�a-Oq�geR**��9~��Y2���H��r�@��w�]5z���W����/.g���N3�e��̑9$�K`��%r��h����[o�&�f2i@��o;�7Pg��#�#��j��L�v1����b����9
z�A����CVS�$H}l�
��Ka/��.�VVs-:rDr�/jn, ����#��C*�F���N�j?ŝ��j���t��{6�N�]�����'�X���F��K*|����%S<��`&Y��h���tF��O���1������F��*���@5� ��i����̼����]��f�'��ݷL/�c(L����G�Y1 ��ԍ5d�>Ӣ`�.Or��y�=zk�8�P�����Zl9-�1nQ�D�D�@�Lʈ���o�~�edg�Vm�~�z�5���*0�c1[�����~Į
5H��A�}� O�{7
ӳ�ubr����+;�^I���X�,886��ڭ��V��Z'���i��?ר�%�yi�q����!(��e�,{�qdGP��Lo�����z�(7p�@�_����̐����z����Q@��i<(�.5����Wo)G-��i���^��At=�ar��@���u�(��EǄgR�nr�x��+=!}~(+�)�DKxBqV�?S�6$얎W��^�*���F���]#.���}|��l�#r+fj���r �q��-�� z��Z��h�}VE�d���"T�M6�gA�3�4���l$���h3���r�B�Əg�����ϩ!>����v �Hw,��p9ud��|k:��ϫΤ�jP,/��t�f9�
+4���X%M�]�",J$D���H���+��}M]�6�ל��o�Ĳa��ۻS��Py�0}ͭ��H��m<p�;p\sbց�a�&��Z5R��#����e��|s����aD�`� �F��`Db�l�L�
/l�M_k^mdm�GW�f�z�=�D�.Oo'E��5�!��P��[g�r��$E~�n>ȸ��5M�
�o���:7�ؐ;rL�dd9�tad����r�ga��qU�=?�R!$J�WbGIl�X�����1��4~OIޢ�F rIY)ֱ��;Α@����	��t�%2%IE��F]%���lጮL3������6�m�Z�s��1�������	mQc�O����W���*��5[fĒ�����Q�9)���j�I�
�Ub;�����:��x��|༕��pVJ�1ɸ9Ufu�KTA5�Q����'j�*���p)Sl4�l���+��So����t�(~�UDu1��^���O��?c}7oUT~x���H��Z���j��%�$v��k�L)ޛc��ʶ"������LA��1����ź�:{Iz����o�f�AK��U�<����K�[OM�540?�ա0(�.ͥz����n2��R��{-�&p��o�8����Լ8qC�;�8�Nus4��Ѻ�}m	���+�����C��2c�#�+�J4�\8��
�x�"NS��f"	5���O��!FI�Y����u����3���%�!��َ?�x�MqI�0��������ϴ�<� �~�`��K���}������$�||�BI����������x�/_զ�bPۗXz����Ө������̨���|{�p�!����/��#��imP�Ԋ���R����xO��t���Fx���������5�H�D�4ߢ�;��q�u����I�fC$>�+�[K͠�Tes
hd�����M�gl:�=C��Yf��'��9����}��]��i����!g�)�!�&\��@�ϠC3̖�dL)��<�ˆ;ٞZ���(�2%��gF\'|`;]Kf�qEx�f��uJru�����Z�G��D!�u��RV8m�d��02�|#:�P�1kܼ��JJ�?�+��G"l�����Xk�k+�[�G/ҩy�1�8 ΅_�/��C�%�̽2a�V�?�ȶ�[6ޫ#me�v`i'5�$ԕ�K��6�]p�b�h>@<���N�׵;�k-,�Dv9\�*�5�Ü�^�znn��_(�i�\�c��j��qD����/q=���TX��������S�I��nR(E�Ե���{1���yS�D. ɽ7v&��m�H��D��*��������H�0,f�®!�����D/�G@F XfI,�'4m��(+���&��.o�vR"��_Ò*]�u���rja�IS��痚\=q��껵�U?ɏQ�{�S�(Ӯ��
j�Ȟub�W�ŀ�<k�ҿZ*�\飺fe��
�6����&�ph`��pm��A#Q�L�uD�s�-R�/T]?"�U�uc�0�v�eoQ!'ϰ&�Ѥ���u%ih ��H5����a�7/g�T�X&�>�Ԇ:���4��y�l���~��,�6�sg�4e%��({�(t�N�G�J�(6���A��H�L2Ka���c,U(�A�=ӿNo��z���A(tj2P���m�����j�M�����2I���F�0��.y<�C�X_)��o�iC���BD)���:	V��)���>w��`X��	��p1�lJ��&/��(��b�Ѩ���hL�g�lC�xo`
�˹̈́�zr�@Ǫ��]�]=�4�)Ƥ\�E<p3e��ʧt�/�&��0<�j���1.�z@�v#���"�u�<O	A��Wcbp�+S��,��wǂ�q�q���ei�� �^��w�L�	?Ι�K2F˟9�q9��Y9s���f~D%g��)ʒ�I��ʉ,�����0���1�,� �6� $*e�^���A�Զ��5��1�ο@�$} ��"���>�q�?� ���CKH̒�*�Ȥ��Sn(�����(��D�Ȋ��d;
}�|���u�Cj?ze�"��L�������D��1��ĄV@�[���<ߞ���o'�[�7��Z��IP��_�L,�ڏ��S���c8,�iRR>�os%9��W#E��ͱJ"������ �w��G�t�Ш6��V��u��H���V%S�ģ��Z���$�l�%�])��aˊ���ޔU����"%�3K��4��@6l	���4h|��޹k�_$ׁ*2Lœg�>3q_�ЁH��_��@�iwP��Vp(<�;9;<2��oN��$gy�T�
T9q#�+���SF-�2�sIRm�3&����&w%Kb�n��P<�3"�P2A��KH���.�J�w�s(ۈ_�'�q�·{t-0�����\������0Y��8;�:K��<�p>k�I�dS��ҤZB �=�5%^p"d����~b�'�^�z��92}-\L�Dp�η��ҫ�&	�U�i���`�h���M�������͚�F�"�>�<�W�x� ?p
l��;y���"gҺ�MX6�j�ȥ!�mT�D>�W��rC�v�}?���/��bf,�	2�W��r-���MXa�G�;�X S;r�J>k�u��c^����[\U_���3�|
W_���y� n[�G�ey(U�'nA�݆#��?E�Ő.t�}8�"��*:�xr�Dev�e0Pj���D���Fn?���9I<�P�g��K�����E�<�����4��e��\ֻ�.���eNg�YQ�&m�=��r���uq����"��쑚�E�S���Q{/����tD�� �y>4\�͵=�,q#�!�A��>����#B���������["�t���ȥe��J#0�Ets@#�����/F�֊B�E����P&���{�OI��UCϹ Ԍ���$_F���e�q��z��ŕ|�Ϗ�GA#G\5��V~��f�H5HAl�'y�-�ݿ�{3D��y���1tU|Z�XC�6�Lfx�(M�o�5���ݾ��H�4!^�͘Z�5,����§ u��#�Vh��fJ�������Z��.ʡ���/P5R�+;��5O,���PG�a"U���çb��<q�_��N��!w#v��a��3��H�jʍP���p�a��&��9�  M.k���ȏ�.gHa𞠖�C�����
Χ�{���Ƅ)Ռ8�jo��gH�����¼���"L�3��#� �M���h��֘����)�@�/�Ƒ�Z.T���tH����v�pk�dԙ�� �)]�ś���z,¥���uC1�Z&�g�7�������Ϗ.I�	,�t�6�ֱ��-�2�HV�7��R+%9������5���)"�`r�%��y�o�qny}��e��h%S'�{��(��Ԩ*��K���TR;TU��ȼ`���V��nNay
zm��d߹CRl���̈́�/��VE	��������JE�-��3���3�&�]�z��=�i�i�d4I�j1Y�����UK�*�!���F&CE@fUp���%����R!��ޞɪ������ ���M��X�E�h�C�ž�筪����m����s"��H����n�P�]a�X��}� U��rӆ�I)��vw(_�RP����'�}�G�y�6��m1TE��6��\��<���wL X3$�Z��,�w95C�\4+�������`!�I���o9���V��Y���e�#�)�ʶ����3ҋ��*�HgP�>F��h�ɓ3n�y*�A�x�34'��£�����e�	�؜��v���OH&2M�W��j9T���d}M,�@$}R���B�in6r���,��f�V�s� �6���o��L1#%�<|�WW�P��DdG*8S���r�KǺ����[M!�9z�;�N�zsV9#+oo�������[��
�� ���U��Uz�Й,��	�|�l�p8�]��a-��������16�K��O7�(�L�2��ĸ���7[KAٽq�'3���>�อ�y��#W}�������p�o���`M��!m	��
��iϟb6����H�19����-;���q�00���'#�w���S���;�x�K� vk�`3PwM�ՈZ�O����S}nnSM���ì�O^�z�l~��U������7 4tե�P{rw�Cv���l��Q�q�aI���qJS �����
zf�u�h��E�I��q7޲\v��%��M�k	V�����S��Q^@��m���Sa:?�qB"4���$��b3�'��-�Q	�J��<){�JH��+9ZG􍄸�p�����<��)yl�O�=U�VGeS�5�&�f<OV�Q��ɑ+f�1�2&�^�Fd�2<�h��Ʊһ�NC�g�3�Xd}� Q��g�S�~ }�+��`ч������+O*���n�J�����I�'�r��j�6���#B�ՙY-N��L�k4_�����seI��6M���a��ߠ$T.|{�>��q���G�z���- ��b$���B(��o��e�d�Md��P�/���Sܴ�yl}��Y5Pz���ʐQ�:ې�߾�E�CcbX�d�l�������av�U-���|�_�QZ���1�m��'�*��5q�DЩS�M���*A#��yA�m�ʫe��REi�/�5�F����x�$<FS�g-k	7M��� ]p�I���f���7��v ��|��C����	͈?jܵ#	�m	{������7\�Zq�0f��Vw�8~��a�|pѮ����zu|�����Q�5�o�ez��D2M����j���*y�WZ^�b�r�z��p�w9ӛ��D�nB`� y���Y�&˸+ ��ǇNČ��R�޽E���z���:�}��?x
DK^������^�A�)�g�����9�~�8�챫M�M_�⁞*�JX��*#���Q�3�i��sX�y���;���ڠ�.~�i�wc�:��\�ʠ���4����y s�ٵ�Z�A9vO��hAM���Á
v��<xyܕO!�����p������EF%-l�K���BA��'�jl4ߗ�D(>��>y%J�%f��#�!�0�n����p�l1^�2NS�T݃� �)�xPS���`�4]�n�u,�+�;�Pw.�<e�
�H��%k���4:<Q�W�zb�$�*p~�j7Z��GU>��y�dYe�8�j�+ �R
�����Dc/�.*>��%eS��a�����n9������$�-�h��r�GIȆ�j������H0�P/���򔷘��IsQ�(�P(�y-��^(�1�[�,q�R��pn�槏����׺�!�L�C��"�����d*#[�)q[աɑ_XM��7���hzA�2i���5�C+�%���B$��[+ {����֘	���w��y�~�>��}����n���
�!�o'�M��}B?�aC?��;����:4��d' �:�h�vr�۞��>T3��66�`�o�*�)VL�I�:���{J�[~�z�h��iZ�]޹vmaE���>C�9��k�""�&���[�ă�nC� ����޲=��,j�ߖ����3'9�����k��F�v7�7�j\�����
(�?g4�⟜�X�������\w�ӕ �3?�F��Mo�E��֚3�,8���E� ���WϺ���k��OY���m�
�ǭ�C
g��}���/�˴��v.���7�[�G���	S:n������܃�F��۴=����h�J9_���W�y�D���U�2ŇQ�7��G�S�q�`Y���ԡi=��-�6c��9���w�(c��ԸU$<�vr�|^l�ػ�G��z(jc:��d��&��KXg<o�k�O�gx}�R!����L�]�+y���#B���&;x){y�ɳi�].��(w�+����K�F�"����	~	#���}=0���X,�H�<&�v?�}�F�&��\�n��F�˂��M�?&�ʬ�l��l!�/�b�2�b�2h�H�N�gӇx\*~61�/P����gj<�Ψs��'I�yA�9(c����5�'Dh�y��|�{��s ����zDc�p��F�$�\�Ю��. �R��8'Qn�8\5G�
�q�y����'f�a�5 ���M�gDO%p|@��.��m�G�qA����-~,�BA����g<'́�[��O'���KI$�a�P��?�?�A�Fc�/��-�U�+*] o�����4K�g��!�P���R����#�Q����g�k
��9��Ph�ו��i�m��ٶ8�"�����=9�+�R�Q��E�	�IfJ>�.���iWnH��9Z��zR�!x��8���\��H���&O�Km_J�f����U�z�����Cu"mf
�n��(=�����FR���9��6پC۲��KN-��^����y�4D�+�tVYTaj� K�Px߰�y��_���Tr��z~�w`[����������&ͭ� -G!3�"��>$��?YqkW����� ��|����{���}��h���I ��)F\�	�6��92�[Y�WZ��Q�_ȼ��=�5'��V�fܳ������&�t+E�'w�ib��	;�D��R��>D¾ɸr�20Jb�r#��>"3"���+��ޘ%���K��/8�Ħ'�
�R����$��7�O�9�b��;Q��)�Ahyz;`��Mx�1A�N���˖p@?�
���������P#��5e��� �Q�H!>�-^/�+���Lؘv�̙����\C���"���}�l?�U���\�_t�[[��&R{��=P᫊��v&�K�h��iѓ}5gR*�7V	n�ֿ�d�m�y�R�Jֿ����=�>�Ó��x<�EW,+3�h�W̋��;�Z|�CQ�.�˓�ft�K�lT���M=b��G�l
�v�ݮl�n�g<U�^��2V�I%=�+|v��Jm���Ѱȡ�(3	P����iۥvX���N��9v�4���Xq.$?�h��sN�as����yf�?)��Z}��`׿� �`#�U��m��,畆�ķ����Jp�0�����ܞ����2qH�j����sC��-y9�H�f��21�}ָ����)��{��X߈3���P!a�.j܌Es��p����F�Xȹ
��N��7�ܓ�&5��0��Q<v�aœ ���k�?���)���@,�&��q�s9jZ0�}�X�w�0�lL��~�ٓ���f'���?�4u�q�C��g�E��т"C"��w(/���B�8�x���w| 
1a�ș��N&�+� �G[y�c����S�Տ���]����q�"�=�P)�&f��o���)vW9���AD3��X�������S��0@��N��N��mq��t�*VC
?:� �?�3�Ȝ��
�����,�6�g���;�ɐ#�S�~'ւ�s���:@|o�e:5���C�"6J��E�B$}����}ڙ^'��&�
����>q hQEP�,G�l���W�"	wd�0����k�*#�dZ]�`��� �X׿��U��(�ijS��d�?��Q�����<�Q�ĩԢ��eDP��L#�-C=gÎ������
S̨-1�<�T�d���D�}@�Z�c+A!X����ך:�0k���٠y#z�4�Y���TtZkU>���(0%YT�?z@$�r��aN{�ە��Kdb�U�G��z}b���}����&qͺ�q�s	R^w�w_S��b{�㽅@�V��ִ�U�"h�k?�w��H�J�v�B�Im�@�7��*�*�U��NQ���`��	�>�x� ��f�M�}�I,�}��0�ES]үo{������������U.r�1?���B:���"�b����[��d#�b`��|*���r�o�.P�\M�|b����Ƞ��8�0��S��N�%�n���_�IA�)CؿnUf��=��j�BXN壥������o�-6��Yu��n{\��4���{b�}��	<O�VLSG�~Ť�&��}���4
�b_0��&�E8�%�ԑ��3EgoNx1y�=r�,(P!��¶���s�-7A�f>0n$�m&I��4,X�3����W���(I�U���'��T&�����XY��M�.���e����oSo�)�oٔ ���8�7`���cK4&�M��}�O���E����B ƾYEPI�y�!��t�Ozx�=k��[ś啻��ƾ��f�����v�@um1��P2'��g�1�tKQ�V�M��f�3[�?��w�l�>�h���� m�8/��z貋w_Ą�x��0_����vő���7���@u�����O���[�F��ݾX����r�w����kIj���� �\T
4�/�������bq&�;&<�&�"�|�Xy���Vl/*�g�C�W����$��K�$t��m�d�HȨ�o�~O��{�8�%3^�ޗ.�y�ӱ|�}?��o-Su�/A|�~�
tה�[oL=T���dZ������O�/�����?B3�����ǅ�B�R����J�~��o�8���%�A�c<��F�8
	(��W��D*~��u4����XA-A/�b7$J��/��wU��峁k�uI��Z��M�e��f?�k�U��l�π���jq�|i����������>��.G��j��y�E���N���!3Nl`���`F�@����ù�#C��x��}��	@��A�F���0c�m�3�(��A,���Fj�P�����4�N��5��ʵx��-����  �:�PO����͆���(�o��ocM���n�}��X}�}�[7�Y�Up�����~ ��Nߞ�Z�Ң���s�u+�8������J�9��/J����_@��� ��J����9Ԣ��� 6g����QqX���gIFP�NZ31j��������8�N�������֗�k����Aa��Nx����n@�����N�a��0��<9���0n�8�P~=т��5y,�FO�%�q�qzCs���s���e�Ôp�MC[h��vx �5]���2��6��3
��Ug�zo=߂� Ļ�ڌ��N�ڬ��4�p�C�G�H��l���C/�0Ow
�"��-����`�����&m��ln�����/P�E��y�s[Z�C�����瀔�-�k��>2���8}Q��ף���>�p:�UU)�1�O�n�\BNV*~���<U�ɕ��%	�7�� ������EjZI��O��^mX����n��Fhh�9��c{4��8�=n*)�K�8�� �=���t�:��X݀��]W���H�P�de8��ڞ���᛾�2���t�#��O>����'*�o��r�'%�ԙr��Ir9�B� ,&;��]~$��xt:z�{�{K��Y�G��U���A`����ީ�kp�01�@fO��<�]W�3����V~��> ��{z�����˩3�n���dI�R�d��8���99ԍ��+�~�ע�&�Tէ@qWJX�ˮ���}$�ڻ9'Og^��X:�O��,u�Tn\�S�!ru�0���b5��Ʃ�rǈ�P���x%��~+��5��&��L����v��NE�r[n�Eݎy��I�ZFD�Um���R��ϩ�|�)T�c�%�����bM��s��%�T��Ȝe�����!��kxt�Q����w<����
��.�jƝ���o�o�1�vJkxeȶ����ai�
5jX߽8�����X���a&j�n���f��4��
�qzXz�d�<���T�qv��kX~�LzvG�u�	�6�SD��Ⱥ+��:�]&[�{�-�{x�|[&���x�24�������O�z@�&�Ҩ��'/��1�L���7��do"X�"o��>r)$��.�U+�n�_t�S�����0����W7��=�����d�B3L�R��sv��dS�O*�j*���8l:�z'� U�K��P��ngG�Ũ������i��yr�\l��t�E���R-U^֏��Q���j�-�����k�2�8�|�4r��p�V�!�=��-��f�=g|{U|K�2i�71��=RyZ�3V��Sj��W��[1J+_@�<��Չ|�����-��3A:���H��H�(�ȵ�Ͼ���:�����`�^�W�wg��	K�
�	i��0Ha�%��x��ڊ@��k�2l�c �0#�#9�0vt��~�T�  �4��6S�tҞ{�7��?����w7"�j=�,֡S��	^B�tU�֣Z���qX�*��>�*:�z�5YX���͞�r��,�&���S���m��8��%Y�����N�������Ԡ#S}�r1�P���bh�������� 4�t�A[� ث�0-�	��r0��&�Siw���Z��qK�X>���A*)�ad}�*g��O_�"�c�7�`1jl��G�þ֨V�Y�'�e���k�$Ұ�i��Al�}�nKV� ��9Z�(IP�6J�%2=ӔЁZ����[�"jS��O����kG������`��)\�	v���k3jt>zE1��DKn|�RMD�0���E�Z���i�qb���w��0|ex�#�dM)]��Iz?;��N�P^�b_9�� ��h:�%[ji(A��I9�1ؖZCܦ�Ω��lA��z�{Ԯ��8.�݃����i��$��¡��~�?3�ki��{��Jњƛ����/ĩ�NV2�=E)Y1� ,3�U�@��AD<M����6+[Nʬ��'nc�ŚE���hN�iL����*�n�r�;�;LL${l���2��%��u]G	D_�aj΢\�aj��vDM�^^�M�E�v^ҝ���x
����P�`j��G��C�ɻ�z�y����+���2���+���U��e��V�)�<�إH^`�t����i�0���A���=fo��^��ߑ�oF;�|:��``�M�j8������O�B��m:��E�(W����M96�R)�d��~�0�z���A�JQ?��������Ư��큺�	�����,�i���L?���6��VlS`�"&�}���&=4d��,o{��}vm1d�1���
W�e���K�s�w�d2��˂�Vh�^%���	��O�c�������9��Z~NW�� �}ʿ�p��RV�gM���.�tX��@/ӮֻA4 ��H�K_|鈏�\�
�{d�$ӟć�J�{�}톅��Z%���&��&�C�6iv��T�i��>I�6�$Bm,�n��:���X	#�a�0��-|��>ēd��C�]V��J"�V��*r�C�*5�:s��q�H��k\�6d	|�v��÷)͇jZѺ�@r�GO���S��u��������D���7O�+����7��
)ə��8��z�z�?��]o�p�VqE����]�s�`K1\��|,6|Ȍ�fEp��Aʉ����"r�_ަ��_�=>Cs� �S��(��_�xe�+P�b���l�2�B��33�9�k��#i6��Ys�#7�7�{.R�ӳ�i�~���o��JML�?Ɍ�|rb-7▙�d ~�Q����,�75s�J"W��Y��E�Ύ\�p4o���W&�P
���A�۲ᓚέ�k��B�L���w�'�2��Zے@o>�5�4�tt/��p(���|Y}6#�3im0`����SN��r֢��r��q���N�Z3�rvR�$bk����n�c��U �|elgv=Qf��/��T�]�����!��32������'���w~�w-��A�s�S�����}紒y����?��^��A"JɃ�
2Zt�?'�A��¡Όr� b����l4����3K3a�H-k2�߻�5�{Ri�m��J`ץ�Lc�Ѵ������R��.����P���f���?��m��jwu���-@F S�ȟ%��ԅ�yS��.�
�fs]N~-�L5�a�֖��8�/��R�6Sߗ�m��[�ۗ���k��t<�� Ȭ#����#۝�#5��V�o��>gA�C��w�z�.bs���0R�T��*.x��*mjLZsb���U�C�UN,i�!�B��s����Y�%{�T����D�Pz�vQ���
2���]��U�Z2���Ȉ�y�hY��B���(F/��-O�+�cބϩk�@��-���W%1?: ��k����D��?�Zi_%G�[5%B��	���VPF��`J��X��������2����#s�Jy�Y~LK-��0��{m� �Q���GQ�Ty�|�Z�&{��<�h���ԓ�C��<fKcujR�z�.B}%VY[��M���(��gM�((��"GN��:i"��M4���@ ���+�����Z�M���cK��꣔v�_�F�UZ���g/V�e�į��L�K�B�)��������>�f>��]��|���?+���x����s5��\�&����"�u�]4�6���;܎þ�6�$ʤ��;��{+^r$�8j�j�}���&��[)!��[�^� o�F���R��dlc%a����ز�6XL�y�X,6g�J������טdAU!��^N�|�� �[�o}{�k\�	U�O��Z204B�SHOVu���	(�^�#9;�c��H�B]�?�D��Q�ҧ�G�\��b�,��7�`p��ҥi��R�����G�g=SVD|̇�ߏ��%���_\b��4��g�U:(�C̭���r,D�(gZ��?�ޛL�C��<�\��gI=A��]XU�N�(� �_l���F�����/�z	�o�1O�_��J��>ϸMgZ2�y�C���Q&����ω���	O�I��@�ԁ��U��X�ڍY�-���U��=S�m#=Ipg
� Q�����1z��/�@L8�+$�#)��;m�H�EC8=>�!�+�93:7���!a-�!� )sǮ24��{���5��b��M���B����K�L�a;�G1�N�;�r���@Ƃ���fzX��<���v^�]��1���Yf\�b� ����N���@H`��qZ�r�2y��Tc���s���,<~y�n��mvԈi*�]A�����l�>}�n�.i�4R:;܅J�HՉݢϨ�鵐����ghƤ�Q�_�7hQd�
R�4�)��c��נ� �&�S�	����ְ0��m˧�K���M�&��O宐���q(>jMw�SM�-��12#�7����8��z�,r�P.z�vpL��n����*�!o�(1k����i������h6ʓ��*-mkwg(�w_��<H�A�#�S�Z�}Y��oS�֐� �_��L���D�š�%��w��1�=dvnzt�|F��Zo|m�'0Tl`��iaQ'�����<̅x���l�t�:����~��^.���%x���j��l}�/�=o�Jo���c�z%ѴW�E�/��g�
}7rT�S �X�[�jn�� �`�����)2$~��c��L,�B��[�����3^��v���S�ؾ��ʟ��Q�xMd�b�j�3��a`��i�}	��X(�9��g� |��K���_�5�+)Km{��s��j�?�zzx��c,�G�(K<��0?qj�(�w��~c�ǆR����s�r<�����v�:zy���o�"�V=
�x���8������1% ,[�Uc��H�Uo ��1Dyz{��.�9�Tn�N���!ג� @�L�#q�ҥ����ң�(0���B▪�>��x8���`M�CZy��S�n�BU>�ͮ٪�WPLa폻\UMڼ ?2��%�q��x�S��|�Wb�Ѣ�u��:+�i߅i�[0�+��7cm˃���؋+3��»,���KDx5�wC^l�Ea7)֦��TG�!���M�Wu��;��>%�"U@�X������7.:�\��=��P������kdQ��!�>=a��m	�d@��)�R��x�`\r޶�E!ǚ�C�$����c�ӷ�ť��%�sO,��Nk�c�J�=����1�Y�r]p�+n�����G��aDJL�S[qr��dZN/{|}~Q�U���R9���%׳���"q��9���G�͈�}��N�����J?�"ߴ�{�����6�����ۖLwvm�������N�đ7���2sH�`��oWEl]bH9>{�Q�Fķ[z,#f��_�h�^}�� ��zt�)��a���";s��M1�S� Uz��jȶ���h:�{��@�X���p}z,�{��-IڣGbg�$���נ��t�5 �ȳ&���2�Q�Ț�T#5;�P��fM�,�%MR�&����/�naJ� J@��ت?�O^�,���jL�WQ�x��
��o���d
E=E�-�C��;�`�?@J�8�5?/ԝ��ov�-�;A�n{�a4Z+t�en-�(�x�s�a� P�**�k�ޱ�Ql��YЦXA�|�_�e��5^�%/o(�%��ڭ=�GM��N/�^G�������`��@odU;pK���e�e����(�_h����wqhN��/t���ܽ',�Rw�*=���U{��A|�Z�� P<	�߭M���<+��AS#�c�z�1�����1��Jg��|ߔ�EwL��\�&�pI�x�*3�%;�Xv]���pEZ�M�L<�o���������}��h�U`G|k��F22	t�)����P��a���_@�I���s)?��F�ӑ�f$v�������6���k*��e����j~7�� *��)9��7CZ�h����)�]������O4@���V����F�m g�f��$��z&�m�Z��m��D����B�h4�sݡe�SF8+�\"�u64ӱp׬=���k(��?K������/��0�]��wF���1	�9�����ZY�g���ǊJ��ԁK���� yE�"�5���u	��X~�;�F��>����$=<�~�.�Vb"�e�G&F��vm����|�2��>-���NT���"��7gq�5��e6?����#З[��P(�%ђa�$O�K��3ر�M���J���1W��ݜ;����s��)��ڲ6��z��ِi���n+E���x��c�!D%�=e��q�3��9�1�oB�XA����9�lz����U�A�3����%$��@�	~,�^M�܍V��E
�G�1��m��N���I�{;��Iq����:_,:%V���R��;���m����w�A|�Z�y�����:j`�ʴ�M7�T������<�C�-w)X��R8V#���Ѻ���)���{�#ڶ��ۢf�X�[
����!pB:(�n/���a�+,p�$��������VL�)'��=��g�z������q�o�Fs�OPE���Onl�)"�J� u�~����O���s'R��ŖY���؝�'���}�%�|��W�� �\����q�*�� nW�ZB*��P�N!e���,x�Ф�0Ś�l*�d�\�x�,�C͞SG��m���@c��k��z<��d��VݘTՙ�c>o6��ʦ��!.�ؙ����;&Q�Q^t$��y"�T��R���V�$F��T�灃_^7�a'6v���%p+�~��u�!�3#�]�+����_=��W��Gj�H���10����JZ'˽3�K�
��q�h��y;aWL+_g��\�"K`��d1�?�-~q��y{W1��#���D��ۣ�y��r�	��Y`��l���G��M����1��.�NS>������( ?-��$_�Z{������[��Q�%�\�aU<��q��Dt�9�����c�������Q�G�Z�b��p�:�a��c�����Tu���ꍘ��:�,K�u��s��OC�rz^���~�D���A���X���J�\���T�!�@�D)�Lc�D.��>\�X�Ƴ���[��rLZ(�zOF���JG�f���?�&[��z��ԑ$�a)C�]��Z�\]�N�i�/���U����-��Փ��[�q3:kD�I��	�>6i3�XUN��D2�t�ӗI®$\$ئ�����]�R�3C�k���n$�w)]p���y-���\Sm!�K}[xy[���P��,�������#d
�E��b�	i��NgLD:�mo�`q���j��_{��uqg�:��{A6���C�Ը�����X8�+m7� �,s��_�V�(�����$�'��rP|N4�-����z��y�(ҢC��&�ߩ�-q�q�nH��N��Z	�"A�ߗ@Z�56��Z��٢��_�2����q���t��`f�UN@a�M�y:�3���d�Jk��z3��?�rھ7>+gf��x-q���K�|[Ku������B�ؔ�L��5����SB�.�[�K(�p_�Q���	���iZ�����[F�ǰz+��{�����R������Y'f)+65�(-5Ȕw Ќ���ꂦ�z�F0x���Ȯ����z�xK)���������N uY�#��G3�{�i�w|�	E�'rY�Q��&,�&��|~L�k�#�}d��r��
K4�ա��(Gt��&�1��)FB�B1̈́f$�.�_BW�1'm�3ɇw�Vg��"��[ex�+V��r��rҭf�a��&p��(ճ�SlwMPQ6a�� �}�Ow�x�b��
�}�9��0�5fL���E�%�;[n�ť�A]��U��6	kB��n�2��.���>���G5a�T��b��|'�bt"����YHǳn��p,�q�b�i��љ�|g��^4�f�Cc��8O�rE��M,Ӯ�>	N<������B��;r�H���;���AY;�h������NӁ�fʎ����p�r_5n���Ւ3P��%}��Fc�����	� ���bvQ�;���sc:ן���ا��2��;rE��n�#!�Դ����9�"`y�Ap�B�D�Z�*�t���{zX��8I�J��������,�3��϶�Uz�&��w�?�J�����I87�}�v*�� ��*٭��6H��q��P�\ ˩���)�KO{]�������;����.�u�G�3�6�x N���gb���Cܑ~G�M������>r8����]7uF�O9*1�q}� 7���^o�J��"H:�<F�m�`Ȝ��ʳ0Ѣ��H��X�A�����Uk^¥�x�3~:�,>�B��1�	���z��և8iÕ	m�B���`����Ol�uwLi�z7�1�?)iVY�b]ȑ�ԊJ��|���+�����18�tR�5��i^4Z���Kh闘�2�����b���	�:t`��E�0Xo�dweS�;8Fan�p�Ĉ	�Եw���Av:��M��9�#�Pd��rZ����λ����TZ"���v�D���4�frl8U�/S��.'��������)A��7����
�+�l��cKF�*ow�Gs2n��b���P<�R	,`�b���g�M"8�W�g��0�M{�.�N�1�B���^�!��Ӟ�/�{t�Sd0�i����G���fl=�쟛&��I�;(x[o��@�����o�m�+����jk��p���$����z�5<B7�R� R�`�*�I�%�a�Z���{5�q���y�#��z  �˞K�@�G�>�pM�,'�X���ͤ��F��"lKMf�r�a����G3���
ꫴ��4���δ�+֔��ߵd��=�>�6Mț̍�y���0#9�Ӈכ��I��O��V~�'��!�V�A��_:݋�h�R\��	��Pz�v
�G�9i�3��Qi���Ycǭ�}���;Nfܓ��[s u����5I�
a�|��3?C(ˏX��$�ۉ���	��z��19�C�Rx�x�Tֳ&��4�U�X"��!�izYM8>��)�#+�a���\��6��&�yn5�I+�Ά�����vJ���F�O���]
���c��Kx��
j������Z&/-�v��X�<��3�6��3�ֱpc�nK�����m;�:���h^�JY�ghg鏷�[BP}�Q_t��q�P*-�-oߥ�}�����-�::%�p��l��P���ߤ����Y�W!g0�U����,�]NV��`$c�� �izFK�Ѥ.���Q=:��o����+���V�G��IR�z��.����Q`��\��D�T���s/\��1J�)�T`�MFG�nQe�V������f�L���x�[���z��&]Jd*x�5��I�f�M����aY��H������_�$�q���ڡ�;�"�t�ad��g�.Ǭ\�1��/r�0�b\��t'�4������`�x��G�s�<a3Y$(lg�Ս��D�Rv����y��C�����(����a��F,�h���=�/�Zf3dԐ�(>3��;HA#�����|i���>+-IZ3~h1��CR9�ㄠ���,1��_�w(��y�	��Z��V�]-�O��NE�`�-�i2(2��P*k&@ͤ��w��&@f".)�	^9Wf�b�r!n�H*X% ls��'cy������b坨������k�C��]�$����Ƣ�w�fg��b�pR��@ M{���>}�$�A&>L�ݧ�J;eN�_p5�y�=7'r֤�Oe�B�_�u�Q�N����~D�>�j}R��+!;ݣ!P�%��e8$k�4�p +l���7��#���1P�z��Hfsn@�� ���v����2���f�lKZ݅�?vu	�p�x��i���A@c���F�H���1��Y�U�%�9���Jt�y�Ho��������t�*ځ����H��z�I� ���݃���ӕ���J:x���Ԡ\��ԋ{ơ��3� Wٛ�M@q���mW�n��͝|�qz��,'��h:�嵐�W
����V�1e��1~���y�8&�5�2����5���� "lO����c�0Z��ü��ˋ>)��,�Wb��O��M*W�_ƖV�^��D#� I�;\@�3�ڢD�Q=����b��b��p�Ιb��	!�A@O	�]�v9��⦍yah��94��	5�4�߷�2�Hc.�<5����(��b|�9��&��d�ξ�]��P�	
�B:��Z�N�F�ڝ�����׾�Dل��j+�q24��S�),8�C[aҎW����)�|�&�%9���Eҋ1u��X���PZ��u+��=XƂ��)C���-�y��VK�s���\�$���f��xेW*/X�9���#>�w/�AP�� a���
�%
E����P�Y�&I�6kF���4U��}L�p�荟~n���m�86*��z�rF}^U����j�Y�]�5S�4 .=�~�y���d_�q�eU��WH�6)U�� �W����p�g�s�)怬 �CATlkw�_��Y������A�~^�}pօV�f����Dey�oVu.�P���]��GJ(���a�!��q�E�pMup���^zT��g���3�K�-dc���N-ﺰ���ɓ��{��4h�>Ю�}�)��ɯ�H�c8�GGMnk袳|ޣbv�rز�c杭=9�T녇3y�	<�������Ct�UG��'���v�=?���P�GH&����0�iĺ��R~�i=.�3T�"��t�������B������4"^:��|�������vɥAъƚ,ߧ�h�<�.�\�d� ��@S|�܊#_|����Ui�)����>��x�;9iS�`�h+^M���r�K���<���[����y�\�8�](�s�WYg�����D�J�n����@�N�D����@ںA�J"=!�L���:�h���q�@�������;�V�C+�)���o����h�2l�J	<��<����BLZ��O�G}��DClT����2���^��I�|]���^�Ɔ[���c5+�yj@�r?lw��c�j둪����(��-X��p�����SI�}�N��TB���AwCg_αHF�'(	�G��zS늱Z�n���A��7u�e�����i�N��,b
ӄ���:X��ɂ��#-:$�M.M`���Y��r�핀�d39{��s�la���^v�����7d�=��goǁ)rp/��Ia�w;��ΤU_�����mm�o��ؒ�hS�a����jEV\Y�9+�$P���n�����F���!s܊@���)���`M{���)��8��U�����l�XBbl�
?y��\�\-�Ԁ��Ѷ�N3����0�o6��K�S���ĒC� %�De�o%g����k�n�:%������Z�p�V�d����ow��������p�t,-�CA�˯�,5���7N�U���G�Jm�AzK�5�	������F�6�w�R��0�V������oSur�4�e����񷣢�b�C�]o��`Vr�z��d�JQ��v�i~���ŐU����Ц)�N�=g0n���7���wݺr���!j��5�u����*��",���Q95����^�~(YP5�����?E�b?}�d)eΜ���&�����	E���ك��u�]��J���0��kKD��x�Ȅ����!L�B�f�7��2�g#Z�s\�j���I��58�FI�k��4Й%D�%~e�볳���GhGl��Nȏ���p3kr����2��/�V!O'G�-�B�(�i��P�2�~������fh��r�/����e��{l������Y> MG��I:@S5�z��O�!�ϩ��ԢB3 ��4�Y�˕Қ�k�|JI�H"�+vѱ83ڌ'�d����(n�Qg���2�25ȑ�?n�_���?�<�Px�6%m�G����(�.�`	yR��F��4(�Al�L<K�c�1\��>��H]P�#2/Е�n���ĸ����2��s�o/H�ܫ������� �Ay���;5]�G�W�T�� �c�?�5!��v�YԠ���F�<s�E+��W��'기/e�J�Z\��G��e�-�}#��L�S�v�S%�Z�71<��~j���t�����F�#`��X4i6)s���K�~����XT�I�&�NN�1��=�
x��}s�z���g��]W�^}䐠�{0��ܓcŧ���X�����$�oT~�G0��'����p��8y�h=@��J��("���e8�gn�t��}>���ZbX�?� )��2��4���j�	o�rJ�kL�\=��
Y-Arr��>�n�f=ŝ�Wl[��|2�ze8f��l�@X���T湇��p/��T�Eۢ��K}�,w4
*�k)!��x@T�E�B"��۷�o�A����&=7��
tO
��<��r�R�?J��
Cp7V-������f 9�W����-��p:I��Y�Eg��%B4���K@���Q+��Uġ���[�e�'��܆�G(;{xr�* }�B�ٌ�@L����l4���A�� 7V�];���qڦpq榩���l�����E��l�!6� ����/�bZ־�~�,��������� �EQ�\� Q�̊�&�NK���` ���V���OD��-�^��wV��!s��,�Pn��Ş�V�Ds��^q��ա��m�s8�TY������#Io��L׏�����.���,�:]/��%CXQ<i����&.#l��A4VܪC�Q�-.����^�1��͵�����rB�%a�3�&�HcB#�>xYŢ��HS)���?��ڷ�8����f}$rk�	���uZ�n�	aH#<x��W�vC����s�İ��2��Ᲊ�pI��+Zc-�x���Fiԓ�S�:쎴E��M�'���36`�z��t�(�xv��U���,S�X���(���O���m61���L|6f�A_S��&E_s���h��|נ��`i7����u+k�>��T�2|���/mⶋ��q0�0yѨ���^����:����+I�n�MA�ܸP�T�-�>���C%�BS3�yt]3f��&ɍ��W��A�DS$&SO@Z��w��-X�؃�����%�SR´���{�a@O�v�6��X0�d_��PչA
��m�
9v7��ފ�n���%��y4���ik���1�J
��'���b%z���6,_��Z��cٛM`BQ~w��
�$�	c��Q��( c��y�A��d΃���U����z?�ʟU�}a�������6�}1O�q���22��m8Yx��F�l����p:�����KΆ  ��Άkl��5�K�r��M~'�������8��#�c��[�C�<%
�ƻ`&��qa�a5id�D�]*)�'�jB�9:�G^)X�ݕQ���\.��3p��G�mD�I��Y��������k�M.s��h&w�b肄3��+ׇ��hf�oީ6�"�>p���
4ꓬ�h��DCV+^���,��:y2���9_Pq/HF��:(u�TY����A��C)olYf�}�2���;��<�
č�7vTW&([_փ�MItj��2���8"�ww���<#����{-:(�b+4���嘋��2I�/l�|(��I#�i��9/MQZP�T�]l9���|/V��I�H����g�f��TXQ�_�M�I�X�E��w�2e��ᰐ�%��*<4�����q��1М,�5�����C���Y��c@@h�p�ٚ%�<`����@L��>LI7yd��ۮ9PqxN�Y,�וoy�p?C�|��&Ae����Iq�)E�u�W�D������F�q�&-.L�e��.�'�-�.�TO<���k��fu����r�w�f�E���>(�ϊ5�kΆ����$ḅ�]��L��q)j	�Zj�������;s����-N5�f�l�$��pC"��/QXC������e��qQl�����L.��
B`]4���M�Z^�w.y�Z82�ð������X�`4����2�'�S-v���S!�ë��ٱ��n�������x�H���
����y:�as혧���T�X�U�UX�A��n�T�
���a�s?��~9�Q4=����9��si8���&Z�0�����N��B�WQ2�y&님�0Xnۺ�Z@EM�=@�#�qR�~M��G4�D�wk�o U ��i��bN*�+(+�b�m@Rn�B�R/�ߵ�hi4������ȼ��-ho�Y��b�)��z���hy����A��n�"���]	[)�������m6���m�9$�¦*}s�!�Eϔ���AmI㇇��ȕ�f�s�?P@�=ܹ�YPY��(��:���:�"�QҌG͒�-<�����\��53=�V�c,v7���	��D�D�$�`Œ���D�k�UT;J(J��T�z}�A�Q�Ix�#�zk`b��`��������yw��������iï� tc6>C��D?fpi^�:��q�i$H�_�Q���3���E]l���
*�l�+d���;�6S{2��.��)�gJMv�;0-�0A���53�J�M�;Υ5q-]�*G����Zg9�i��ZN���D#��9�v�IA}w��pY$a{-�2>=l$�Vl8%�E�OM���R�`)�d~k�3c?t�%^�0�;����w�:�8�9��7��>!9Ua�;��X�\�u�]��Q6�4� �ۅIҦ,:e�һ}���&J��6y� W�*��UK!�ޖ��T���[�����KͤE1���Vi��w1{Å���u�бߖ�6!�r�̹;��V��@�]r����I)yp�<A����]�ͥ���ꮣ+@NK���3�_E�}�n��Q�?����B�.mU�7�)1p����	kj/�r;>�MI\����DS�=���:����e]s�/�1:0�/B�|K4|�$��4ȍL����:�,d��?mJv��fUk���迅}.��?,�[8뇇9�ν���QHsF�vi���i�[�h<[0�c�$���|3RO�ߠW5�R��ﴸ�H����,A:ڏ���� P�wܢ~��UwnH�\ְ�1�ɫn�B�U+����[�n� 2t2D�M�Qʚ��0ɳ���=iF��Cw�I��m�\@�YY"%${N����X@|.>�0�^�����C�pW��t^~d��T�dp=��_�5�����r�����b��u+Q��0Q�0���t�<ݱRJ<�\����@"��H��|����-��~�u\g��i��/���*�a���VZ�l	n4� 댵8�@�U�Z�d9U�kpO�f��)��ś�NG���jd,Z���;阋���d���
j��إ0�{���/k��k`��s#E���|�
>�����M�R�=���R��U1]J�� N�z���6�Q)���_@����u��q�d��)V�8��V]�W[l2Re}�^dS��)�A��4�c8�3h���.���35g���뷁GűQ����@֥�p.�k.C/�����nm����s@�Q��5��)A�Z�6��\e���Оg�՘��旔��0E\�q���egiO����6�7I����N}��*t��8�zƈa��fP�@��-?�ژl�&��i<�f��$�C��n���Hh9Xa��N��t�T��Jܸ�29Vg�I�g�}��n%wVp� |";kW��W4A�J|�.�?Ӯ�-�p�{x���yvypd�Y����~S�#u`L��8�J������N)2�9�D�Ͳ�WL':[B�.1SFo�7��B�z�V�j!�q�sF�����s�w�v_�o8i�q �%z(2���`0�Z)���)fQ���oա� B���3�&��N�:����"g+aJ���C$�M�}f@�ΪG�6:�na'��oW��h"io���� ��G&���5v��q!IM<a/�
N�����9�yt�;ܶp�M�hG�+P��=_�TU�S#V5�~"��6��[�1��M�gZo6i[\\Qt�3%�N[T��4�{8��\������G�Jg���g�R�����L��C�G�$'����jv�Y��4`�����y��\mP��i	p�tk�m�}S��K�ȕ�\�|�3�T��˻I�H޷����.
*��ujJ�&�����yA:�~���1ܕ�����LiU'}L�'�������E�&3 �(шZ�Ĝ	·G��bG�i��D���U��)�C����ܯbdH� ���0@�]tC��q�)M�uy������_��+���R`(ڼUX�l� ~^�� :��oH�.������E��s��4]���;6�X�L�.�N��P��́ڛU��H��u	�S�=��ͅ!{B��D&���q:�x>�u4ԕk�sJ?�r���@YK��⒫���b�#����@����o^׫6UL՞?\u�ï{�n���Rx˓1�4��o�Ŗ�4��차UBz�������ϗ�.�L{�������:ܒ }r�	��l��(�w���!U��	_�i��Z�B2��)D8�>~��g���'m.q��1�Aj4~��GP��c�hebg��j���=	��<�97��&�j�av���(3j��|�wK[L��הK	H�Cz��f�|R�}�@�?����e�3V�V����n]Ya�5ȝ�d�j����R6����B�hIeu��qϵ��4S���Ȝ��X�D��;
�C�/�ߒ��:����-.�7h���rD_�NG������՟���cP�b��^E?'�0�5iTy�2s�_=疒�}Ev�dtmV���2�wЯg���i��u&:�u����M",��	���	H�����[2���	Ne�j����j���"a'A�B�EE���Z�s1�Ee���;�J3�ؗAǐ ���H� �~%��%+ʓ�v[8�v�+���.���9��Ú9�c�����/JȢ6={q��,`�V��\��r��ʾP�>��w�k���Mg�&�{��]�gFXv��&?���̊Kb� �=VY��D�#��(�%J4�>K���Z�3�����x��%��#�dع.&:(�ts�^ @�̘0���c�/'�p���d�-��;fGl�£Ƽ?A��-�>�l�u��2�����X����!.wF_�{?��gW3㤸�f�)v�أh���x���`�_4� �h �)�\�fo(�����հ �@���9"9� �����z�Z.��홧�>��.h�@3p��g�P�1��.//Ի�y�!:�c��?9b(�������� �#��9[��U ���eK~Y�Y��1p3�!歒$b���=�Vn��������a��jq@����E�Y/) u�������T�4jwӯ$�@�W~Dw`����x��	#X���ΰ�CT�����ʨ�\;���4R�3�,{m�yn9׎��)�Y���j=��m�D;�mU���S|��i��ﴑ!��W�V�ŹF	���E:���������Ů����{aX0���Cʭ|�;t ��R�͜�vi��6����4I�?T�y�V�Iq{�O�@������^8f��zE_�#*�i�ؐ��+��)�</�@���'Vi߁ �J�H��;>Zew�â ��Ri-�a�7��� +�t��{�f��=,{���)吻��4 Z���0��8�F8�r�w�ȫC���/�A�3�:���t�#B����~�x���g�Z��9~�U���p��oJR��"x�"�sz���Gw�(�&�@H�`{�>"�Ԯ�\7�(��c*P�Boo#���#�AT�D�}�/���O9+�X*]��}�p�װ���g�Ԙ[���ݱ���j�#��o{'�{���j��Y�[1X���j���Ln�O��xG��Q���N�{v}�^iL�EO.4�� ,���z���@�S�Ck+]bٛ�,�*ٷO��e�E�i�F�3-��ڊ�#:��Nq,r/Ҝ��撛
%���ƞz��@�\'#<`$�k�{���2oD�o�h��Uqe��.�|N��Y�]����Ӈ6��R�(GAZ:�$3�{�V�m�)�댻J[�I�*����@��=����t�k��0\¢��u�ܭ)��-��Z��_�/��? 	?򗽸(���0����Bq.6�m��҉쑟�.`�� ��-&QuF?��DW�3��������ek���(�C-�D���!	pEM�����T0��)Mˮ�=�b<D�:"�L��q��~�P.����їR���f
�)����.�Z�9��^���l�)<O�1��o��^��2�������_'Pk�+� Y�Q�5�Řb�_�P<l�H��xn�yR�8g�7����&\{�!sV�޼կ/D|v�����п �c�D�ۓՠ)�8���w Z���(b	�`l�+re��^WM��6yO�Uo��'��n#h��d���'�������ah��pyIo���RH:%�����UĈrT�Sg>��]	j�	U3��I�7��;��bA���=��d�{U���r/i��@�q�i;�������&E��}&���x~)$�AtT��Mĩ�ȧ�� �(�b������7hm︛!9�����0�~֒�S��X���l�G�5�>Z���9O��]4�#o���)�7�=����e~���ã���>;K:%�:��,��}t��������W����6�cP��ӕh�[^l5�+���6�ףc�W�%L=O���[�)�LF��ޚ[�@'�����&j�Q/:���XD��
�6�0�̪�������Ÿ�/�n�C�֬�^JϢ�aɘ���f�}����GM�sU�vO��M�VT3zZ�>E	T��[�A��?�DY�ߎt����A-���]^J��V�D���v���:�(�`}4�hX;,�<>ܿ��<-���Ք��N�`r���#္���ؑgD�G�H�a�g�]�d�ԇ�VM�E�&y~��a ��I7F���߈~*):mE�Zto�UZ�9~ZF����s�ExRm�&�Z~zY�(�����W��w��Q�jʜ�C��X^�n`�Oc9����J��X��	�w��a�o�\�
�n9����t 4��+���a#>+ͯ�K��7� n�D���ci��I�xh����X���#���|�]ͤ)��y��+�a���/���E���-Cܭ�����y0v��#6��fq��UK3�P4	�V������<�ш�;�W�j� bT�����`�q��m�T4��Ca��Z�9>ͅ1�Qg�?�I�d�&���df�����Цg���ѪОX����;od���{
��E{�.������Z0.����S��%��P�5��>vw��0�ב:s���X=@)Է=}c���倦<B��@:�i�n ~�����|ӽ_\w�w��i�
c<�-F����JIR,BS>xEm���
A@���E�H�GiHjL�`@�juk6�!6�+�E�k��+)�Q�!�[L^H���2�hI7��4��&�Ҹk��=(����$�g z��	I㊨'�����cg;�w��y��D.V�����H���Bƽd�"��W��a�XX�?BI��*��nu5�/�^}2f"��xa�p+�dj�o+����>���*�N�%���rf ��}dx#��A>���ؘ��4�W�:����n�!4�X̀�1�����V�$;!P�cݶG��Y�^L���G�	�8�RT��_�6��^'�sM����&�g-�9�k^�g{Й��f�j1�ɑ�#����b���)%�
�}���Ӿ��MS���L�7:��'��P��� 𡄅.���_E��J<g��o_U���ܾ�/��mn�}��[����'�S�Ug<���=��5ka?��PV���e��Î|���_�>����&`����_b5"nIOy����e*���e1� 	.�"u�F�j�}'j�§�bm�V���Q�?�,�E��Zë�$hWc�c+6�o�Y����|gc������S��g��f�e⩝V��V��_B��A��Lu��Д�-ZP��k��
æ����ǈ��EO�7U%�܈��Q��}m0N�7�%��n\Q�����$�Fh�%��/+Zh�eh}�>Hlc��6����1ґE�U�6�!�˶b\	&�h�}�@�T�!�3X�	�jH1�v�!$5���B=Y�*�M�A���<����~j_�ׯT��E`����:���4^�0Se�,�p˕�����0k91A���`�UUU,�A�/t�Wr�aĴ��c�u2�H�b�\m�QPt�d�������A�����K����xYSRGGxI������
x�dU��4q�e�a�IS��8 u�8Omj-�z�B�1��?�ȑ?��y�Y���z"��w����*K�"���7s`C�dYg��:�?n�dΠH"^��z���5u��g��Ĕ�Ŧ��+�)3�u[o�}�.������	�e%u��1�P�Q�6n>R`�rBDk�EH�Y�����
���J���)k�D�ut�������*���+1�#`��j�����AW6e�4��۪x ��Ɓ��E�p��������B�\��x�����0��٩�a��rn�حf�q\�@��5���R�WrQ���%/�h�|	
��r6�����-kO䵰�Q�f����$�,�Q���;��%N�$�վa�#��ڒ��K���S�6�Q��ML���薔�;,Y.]|ٓA��AU���Oe�x�Gp���������7�Vc��;;�c$���Y�Xm�p�s���p8	Rװ����s���S`��2�M�$���5<7��յ�I�j��~.d�l���t�ZQC�JJd
b��������SP+`���Y��F�n<r���%����ZG
�an�����؝��6�@��ǩ<1�T�HN�!�A]X\��z�ȡ�똖��)2��y׸��?��L���X��H����˚�܏��[s ޗ��57�i��#�����q']z�2�β#��#<�t���iϊ�U�\B����]�6���l�@Ӫ�l�l���F]ڼ�RW35:K��b�����9~�F?�{j�S#�^&i{���V����������xF�����Ͳ�	!���X����_^�Q��&���w/��M������Ϯ������Ѱ7@V��܄�T�R�����6h�X�j6O�2�������e�z���X8�����a��_C�(t�Mkq5
J��J�ݮ�x^#6=�Z���0�1�bZ���f��n97��ha��e%���G�ޣ0���x�/gnG���~�e>^!p�M[�y�9�rZ�4��Q�*��R5�g�I��������+�}�d���1}S��)[���_$����"�
\�u�)j�p�,���^$�.���9�/}V&:x�Ų�GQ�A3�F����Lq26O��p�)Hc��3/�ꐦ�~���߉=�l
#�ۘ�d�CZE��Zɂjݵ\�H�}%%g�L��
Z����啲�đq~�ysM�gD`��QYl'�'Ct|�ůUX|�,�_�U��/B͝�t���I�m}$�&�+tn�0@C��qȄvc,�Jr`��S]�f	��()rPD�Y|��٣��}����*,k�]\��؅)Z���`��5�+�"ųx<WhZl���8r��{�����B')G.��v���՘3���P�W�w0��Olq�e��ӮKo�"TC���Om��XxH'7ʫ{��~�q���&p2}���ֽ4،%�?p��E�!n�R�\I��+��vL�zsU�&�	��^ҡJ�d<��(^��	�9��{8�GL-X{_PO�GW1�bMi�<�E"e�>+��v�o^b�����sA 7Tϧ��z��5 �%�{}�	�v��Rۧ�	��6���1
H��a���.�o���+��ѷ�+nj`#6�k�x��>���me��Y$"�T
�����z��wY������6��ܴ'&��2��`�v���o�����/�u�܇T^h�c���vg%6+���x0#�J�?�{,E�1L��O">s:~�s�cE�������m>|��'� ]����Q#�7imiD��1ߎ=�Ǹd��t�k��q~3�,'�l�+T�A��ܛ�S>��#�О�Q=5�q2�"�ә*$��/��N2�0Ey���{);=&�?<�1��5a� ���y%Go��כ�w������V�B-��P����i��F�.k������i�� ��.Ҽ��#�9lP��c���4q\=��Z6=��:��JUȃ`p��'P,��9hӍ��(���nаД�\˹�g��C�`����J�VV�/������mlb>����v�7�j���Ʈ�׽�+�0�}8�'���N�[�z�;x*�b����0�Ü��}/e�ʹD}d��Q-Ж���*���pqÖ��Pm����=5�����N?�₝�%���!�/�idDI��<kW�3�n9m��Y��)�s�rK1П��Č�Z"����Ai� E���p�^��|��xtq�����t���k\y���,���=�૕M�#yGZm<A2C�t�w�:�:��������i����'m���l���r�TbPA6�3ժ=�`� P�d���t�YEٮ����H&�3�rf㸶�3 �0zG��$2��3�h[���6=����i�ݖ�nRD��c����"�T��д�#-NR?�U�+�څ���f���n1�i V�y_Z���o�Ox�A��᫪r�{��J�m�=N&�
o��R��BKZ���K2�i���XP�U�|q�=q���>��F��|Uͳ/�&�S�����w7ܻ)G;5�KV]_K�e9/bW�:��O&��7tn�
ٹؚ�n�cq�}�gi�Ò;�ϟ�0jp��Y�b\o�ZHq8�+�(�+v����j�.��5׮���O��bb���+�͊���o����\rA�> '���م90����gw�4�WQ��9�À� ͻ���e�K��c�~�mg��v�|d�V"}4b@���WeׅǾ��Jh���~��*Hݦps���mȸQ��ܚfb�+���O�	���%s[�i3�<Mݓ;��U6��QY�����C2�a�� h��\W����2��ћ%�ǌ�m�;��ȗR�H������D�y�gJm'��D��K������f*��o�kΌ�*�����!�a�Jb�Z=��-1�N*gI�XB�띶L�WR��8��>x��HQ�_$���]pL��N�����ڨ�W�ɥ%�8��{��*>c��Ѩ61�}Y�&;�$"��/I�i�Y �lj�yl6:;��(�*߰���+	^K%�b���8��Y�^���� �1�U�������4�3Aq^��]����P]J(�ݴe�mm%�����܀��Y�x�@��g��g�T�vm(�s=�%"��B�dc	Q.��.U��5e}�g�?#�L��¶~ |�?H�C�ǵ�4�8Ȋ�D��X�a[
��.fMߓ�F�yN�k��p�i�޷ߺ�I��K��PK1�=v�|f,�5���,����1�1��>�9��T������M� yyx��T=��6/QhN�ƍN*JR��"�>D���Qړ��A��[�8��D���473�A������0S��)�_̿��2�˕3�h�Z{���/��ШQy�]���lf�=bR;{�,�iM�T�LL`��1k���8��;q�*=�-��x����Y7Ǹ�b���� �����/TO���w��b��-ˑ�Y�B��ϊ�&��|"GF�-Yܿ���ƋƢgo�)��إ�����	X�����?~=��j�`W��qn�Zq.!6k�T&XQ��w����wi(p��d�>�� l����Ԉ��,���M\�FQ���`�S��hr>�НN��&����6����M�ՕaDmA��6��a%�a�����S�{�D�E��[�[�?>-�,��LѶ�~a?��C�`������e9��v�8���r�:A��S�3��AY�BR����đED��"�	����R<�R)�ޡ�O_�
k��dy��m�q=7�4㸹$W��|����"?�2\������n~�(`eC{+&(�bnU�u�Uj;U���ڞ��Y@L�[Ȗ�z?;wo���E�,W�>H�NZ�\;�&U��9�|8��{�����S�4/��A
k��.��g���F��!GZ��U�-( \��6s���g}}��l�%o(����(�~�zO��1Tf2nk��1AR��S���/���:Kۆ3,��e�j:Ɋ��9�=�O�u�w����H�Z�u��$�p�B���3�\��4oA�wH�c@h⺠���G��턠�ڈ����G��.�%=�MP����5�˱1ݓ�P��� ��4����S����]�*^۽�U�Lm���$J;z���koǆ��kV�9qjy.��PX�"0�k�#��)��k1��V�u.Y��hj�,�J݅�9���3�����>D�?��j6ʬ�G�B#�2Ƨ-�1x���Ө�B+�;U]Ur�|�����|�	�`����Sf��h{��R;:�ny\�u�"W�]k*�M�;��}#�NM$���Bo��A����.ɂ{��M}�Mm�1t �6�*���f�f��
��w׻�ջ� ~���V�]ҤH\�M6����C5�"���,� h�?a�%/'��	3�@T�3��0�n'�_� ����'b�H	&E���t4�S�H~�)�Եf%�T��b�� W2-i�^GRקK�|I�Q��/�~��r�� ?�`�����_5"��|�/%��+���h��;�O*ZB��f�^�(Ozl����ڈ���`�z�ܗz����'�h�qppU�HMi�����BQ'Gmd���.JH���"P�a�S�*�T:��?��ü0R��[3;�S���^GJo8�!�cu.���nu�� �\�g&! �����T��DF.���aF��t��
��Ο�ʵa�8<�' ��!�&�������iC�gW /�Is��� �o�B� ����K�o�+���+�" �X�������&�q�
�&�V:��&�~�%�
0��KqjU� D��D��\p���GA�̑���NF�2`���X�|����ln�h�ì��Xk�ߠ�r�y�2���QJ�
��Y�ߛ�GEY6��� �Z�T����0R��'K�S��s2�ϲfj'rw�y���^:�ia�v��32��0�3�e.S�p!�ϥ���a#���tT�c��T�3���*�L����@�ޫ�݌ �Z��V�Rת��q��X�Do���lY@w���v�g�)
�n����H�ֹʅi�+��lo�J?�!���t��ϟ)4��΄x�ᱧ`b�Dԟ���*��>7(�Kg���8%�uEmلe���`D�V{]���ڒ����o)~��`� �T�/FMj|6��]��ê4<�>��æQ�����g?=vm���*����Y࿱�Oc	�o�U�s�m��Y�@��Ϋ��Lg�Q�vPFAp�U�8��؉�T  ���5oEJF';�>����]�AtF,Qʙ��
�`�p/�厸uңX
�GW�=s��K���44#�oM:E ��6o[����J�1�mz���.�7�-:�P�I���t�R9�D��?�p&��|��^h�a�{(�_�xR�5yt�~�b�NL 8��2�#HI�a��):jo�o��-cA���H�T6��{����|���lRm��K&t\uW���?$N���`n.���.<~lG �uI�R���z��-���������H>��]�y��&AU����FѰ
��:��ӺSOC�(:D��\OW�,>�~?y��n�~PiW�ő���Hx�"�V��1�|�/?BL���a�������?�u��'��&��n^{�*u}Nowm��$��0��[����N�Nù���D��0;�F��q��NDv^�	��Rt�F�3?�������=�u?����\����_�'p��÷QS�z�Ə�cLx��q��\�B��*`��>
���r�5��p�����J�2.�|ڠ�$��9�D�e�0�u��|Q�'1'V�ԣ<��b�$������^�b�����N��������5a������$H�1�x{n�h�5�N�V!�E��F�D_��q��f�Ja)�Q{a��T�iE+�p�#�k�
����ht���V�գ". ?����K[>PzZc}�E���ht�a�C�������bA-�4���o?�1U�K�����������SL�_��)]&�#���`�d���Ƃ�'	��^�5�XG�^G���m�ߜ���Zuk��`����O#`������'���o�;hm�STa�Ge��$XE���%Z�w�~Ej�k�+�w=�;;�N�I͕?_�a�ܕh:^������w�d��&��F%^�H]`�.A��W��f�pG�9���B�_K���C�Q���9��"�w���aC`�N��l�@і�og��#ݱ3h�)�V�3CJ<ú2|�;=��O�)�����V_�OI1y%	�Jȸ6�IQ2�#*���i$�/3������R�²&�n�t�%��(�-��Z���m�i�	��[7zΖ�� Ж�x�f�xu��#!c-]t�!��V��'h�,��* ;W�X�����
��\2���S��WMI��8R�@�!��Wϑm]�D��>I���0 |��MD�����Jc3�bկ�L��f��C���[L�4c�����H2]��y0�"��v�d�,ԯ�78Ez�32��˖6�>PW: N�ph���R��AI�M�xP�WA䏤@����˾H��C߸����lN	^2$7�B;2���6�c���Oq��>�j��F�i#���yp$�����< ,�e�:6)\A�E�3�u?K�U;��h}%g���v��\KE��O;x��G�i
�K���K�O��zo8lrM����ş��$G\�ϭڲFZNx*�mS����gr�h�+�v����s�e��IOP�f/��]��du�G��x��K�q�@�GI��Y6m5�&�~��7�W8mÅkx��������.`�9�Y�t(�$Y楛�_���WR�܏Q��)5Ժ�����.������Q
ZȦs�[k)�;Έ�!Z��a�5Amr�Z�`k���_I�
�ݞC��#�m�����?�XI�W�ӎ?R2�-V#������6E�|2��g��r��I4��.��LU�V_~S8����Ťx�.s|����@��;�`q2�X���jo]��xP𴢹:���.c�;�i�q�h.};/��f��I��0>����AY�� [a���B���6mȰ�7��J�4�y?��U0��V�cT'�Ư�7�,E]]-\���l
�������xxho�Y����I��ɓ�VZ۱�A���N�w��χ����#>����m�P�L*+��J(E�J�8$��0�3A)�T\k�2_���"z�yϐ�FՅ܋Ǫ���̃�� #d b�wIK����`�g�s�hs�Y�5Š~`|��{Iɩ���b#��`L����zQ_$�Gq��O��n�|�Z:Ujv6b�^����_�*c֍f��'�*�|v��ȬRMKV!�n��b�l�Д乣����J�A��'GIt�A�+P� ���壌���S�������sr���QĳW���ظ���ou'P��/P�,�_����6��<�6��9g
v>��C`�#
����G7]�|�8���0�YZQb�~#D&����Y�$����$�7�wW���4��֯	�|��:Sɝj)ya�����i�~iu#�l��-7�P$J�*#?�_�֔Ӭ�nz��@)l��O�������]Gg����z�һ7�'���AEd�i�ې6(����v��Ae����)�?��7�u
��5�4q�"]H���}���q����W��_��{PN��w;�0/b͛he�ԙjy��2�C��F��eU�V�u�f��!�\�tˏ��g�n�	_(_Z 2��G��aʋ0v3�"�NE�y�p)ǡ���Q����bͫ�t�IF�*K1ԣ���ȥO��A���"��L��S �=�p6�\s�z�u6��Ş�5�W<7$TzzXXY�u���x���G*�mǾ� �;�l�j���К�q���/�m=�>o�[��I��d����� ��1g��"(����$r�(m�u��EjA�<���ɡ��ҽtB�X!k1m3 ��s�޳����?�	$U�b@���A������>�VEc�a#���QַͲ�&�c�b�1H���VpX���q఩��1�A�� ?U�/���L�P����D��ߔ9��8j��%���u������Y���A��vBԨV����k�gf����	��z5rY��e��ƻ� �;���vo�%	8�2�oL�����q��&�H���N�#&�S�i~%�<T�z�Q�+as2����6��z[�> �o�|q^���9���(����:d�����h��xO���wSc4��F'/ ����2�J�Y��[دN6���(B���oj��]�_0��C�F��*h7��}���n�4w����
��5 �������Ā�bs9
�0�T��2s�0]@5�ȃq��,n*6�c� B��ͷ��t3k-8b�}\!���W�e>䦠 �/���m�BԱQ����v}�N��P����^�"ގS$5s��jj<�����l�,y�s�6Eb4<ڜ�����˿55|���t ��fH�/�5���n�bb�!κ��ꒅ��w��3Q��"[���('2���<�����%��Xy A�6KB'������b��ޓ���ܬ;����ܦ��_Ƥ�;E��,�4c�Z2A�� N�	`-��0�+�npn��S=D`P�$�W��R�.M*^�«�U-�Mf�Ҹ�s��J�q�T^�+#5$��HW�H�w�k��z�ſ��ѫ_|�辬C�M��A����O��]���*��7�؈�GI_�>����i�d��%߳k�EӒ�����t72�2�	�^ŷH{El����X���B�R�f�F@��r؇
	��0���)��6�f��poW�C��HݹA�1���(CK��t�fa��������xWֆ:�60E~���.X�N��H3����e�����~'�5 ,��SSaxApE��?���&)����hȈ�,��0
�&��21	͝Cb!�� e�^���������	���(-�o"��Wg9efj�����!���ق�%��0��:M��UC�>zT���<B�[If����@fu_t=e�k|d*mF�X���/��fJ3�qtE�%��Q?4�;e#�`�)������1.5�l��ʀR�z���{���]�b�$�L=-#͵�!�;��L�ד���L�1]�K�U�(�UM��r�q�����[���B�sBR��Ca�
��g�|�_e��Dd�<��w��SEbU��0r}��`� ��kK?E�쀋��P�e4T���xsGѧ��\��,Xs�p%�ǲ��T�_��D�J�`QL�,I��`_�ۻ�h�p�pc\oTI�⯝S�5p�q���"�
Ϙ�6?X<V�ܨ���F�@�5��9�k~d����S�>��'k�#Tg04rAO�=i�ڿ�qz��K\տq�"�zMo��Q�; ����eK�1yBjK��j�Jq�1�^e&x�bK�;��&���g�s$8�����$�l�(��#c��]��H��'b��������@��XVb�L��{�i���������o�lz� ���Y0t˲��s[Gl�+,�� �G�;�~¿Bj>3¡ǆ�6��t�ZX�]�kL`�{���ݶ#�\�v���#AϘ�R��B�k�Ʌ����怟tVl�T�������c�]7�p�z>���M۷�$��Q~'�6���_�^`�0u��<��j��Ě: ���=\��h���6�}�K�8�1�t_Q�l�SDFG�"ŕ8��U/�Mu�$8��ɷ��c.�a��HKn >/��y(6���=	1]�jV��t�+ �P�k��)�J}��Z�F)o�I�m�MI��Ѝ-)��ʆ%�LY��ͮ�x���CH�晘��Z��r /�+�u��n��Ow~ǹ�mp��}VZ�����
��d�m�'�E���	�M"b7;��M	 l(���^�)��o����T��G��\�Cq��N�­ůF���Ww()�Mx�|�P��v�l "4��� e�Qk�c�A�3!ґe���"_>�wh����C����+?_6�,��q'��O!��Xa�'� 
��uȧ�Q]\^�.|$!F�
�j!����BK,��`�^pZF͍U���������po����Qf_�#�zk^Bq���\H�oX�B��%0���J�ޯʷ���m`!K&yNU�1UD%Z���^w����9dh��u�{���f!���_��V8�7KwMvD�H���-��X�n�q��f�Q@��Vd=�C��h���_��~d����:��w��Ȑ�]Z�eil�'0'�[��e��,.-��
#>�:�e3@��� �VX3�����cK����`7�AbRF�N�����ŬI�y�F��M���Q����e�#�&�˻�䷉k�P�6���G�������]}�3�h�<���?�c
(�0��IS�j9v�:�X-�m��̫���Xԑ�M\��b0�\W�l��-�^)�t_y�.�&���\����;�i�B|����Lb�Ӭ�C"[��q9Lc���K��!�!2.k�����]�Lr����U��J�(Seqa.��VR��ADD���&��!��O�L�/2��۫�Pn�H R&��r������RF�rA-���>�,�L ����-�[a��1E���Ŋ�^�I`g��T#�S�z&+ƥ���t�@t���Y,V��',0���j��(�'P��~�L]��,;�`��*hx��8���a= �E�zX��;G#a� ǖa����2�М�2}������8����75Y��:d5	\g�dǆ4'>��b���6ȷ%P���`�xk7�2�ڏC�9O�I��g���^2跑~��[��>i1;�8YA�~#Ů�]��N����ƯTys�F�_}]{���Dވ@V��x��TG��,w�ɏ��@���y%"K1�Ӽ���(p���؜^��c��Է��!���	�0K�i��b������b�LT�˃�����e�%GF��'p�{��9�R�U{��lx��$m.-�(Gªf!>�컒P���^XB26,��Q�:V$g	������^��?��cb ?�=����{
 -c�6c��|s�R�=*r��zi3�m�l8w僯V�������q�7����Mc�����dǇ�r��ź���	���V��z8�'휬�����;��E�a�W�mY�w+�F�m|8<{��>�|�ч�S��'F��� �.�l�2��f.CD+xh�f���>����	ow�yɪ�IX���|U�^s�C�E<A2���#�w�!*w��z~7��Mz��_.�5��K�x��`�M��4˘���c�JQ�r�Cف��o��^�/`���]*�1(�!��k"H-��q�c��6�a��sۄ��������Aہ��[�W��!
�@�p��+�.a�����B�n	�)������<��k���6n7�h^����H�ȼ<�҃�((��[��TF[�ԙ���C$��X�zL�00G@L������4�ݢ��8��d;M�8�.�w�#����
�@Y������J*�սo?�C���+8�h�9Ʈ��FA�9ө��n����U����w����1�;�%��ABIr7I8�_W#QD�v?�Euv ]rرF���l[
$��U:��e����c�i4�?�	�U�Hz}+k�c.�q�����>'�M��ՙĵg��ú��9Vz5�&H�K�M�k��:^5=27i� ����Q�� �G��=ҧh5�՚�E�().!���f���0�ΩG��Ì(�\-���#6ߏQ0Dݝښ�����|�sq/+����ҋr�`���/��뷯ɢ�h�� :x���S�c�[��asL��BD�IV�X��\y�k5X�s�{�
�.=\�I�O��I���v�<i��'�[�[Y'}��o��Z�i B�*ُxua�{V��Q���F�����Y�וM�κs�q��6�Í�v����@��j�M��\�
B�!ĩ*^̨V�9^#0�I_7��GR>�H@em/L��� %j�S��pv�ă ]c/j|�S���_[����0�c��@{���og�*h�D�`0�����d��f�}x�Yz�x�zp����u���?�q,Y=�jM3��&��*�&+*�8�ϫ��(!T�_Gb4G:�Q	����%G�ެ�,� ����ð�������W`�Q۶{P�HR�����W6��W[�!a��6��vx.�=�F^�7����q���1:>�<XI�*�s{��{n<�.CM�xnvxy�^d1Z�����R�z���L��G��
�+�h���!tcۓ�Д�eod���Ε��{��g��F䗉�_`?�x��x�cy��^V���ڨLd^�r3���&���{��(���~�f|I| B����Ȁǹ�:�H�9�3�ٴ}�J*AhP�& ���^8D�M�ͩf����A�S�t�v���X/�9>��J�4�׆����I�xi �je�ٶJ�+ˠ%j %1��9$��a�.�J�0/Ը��2���U��(Ez͚��$�/��o���ZN�4\k�� Ew=�� �t�`O�qb��E�ys���\w 9fR�����ٔ���}����p�6��B7XG�[f��2�J����7���A���5� |bV3�G�V��7��:zP^��*U�\���
z�'��gF���r(S��lE8W
�{��7:��(����#�j�h��u�x��ch�'N�젴J7��&z8���ɥJ�Ⱥ�IGa�r"�&�o��6�)9|*x�P7IA���r��Bx6��ޡE�D��3$�]v�}\��
�<2�2ޙ��dls���{7E�*X��uo�q5Ъ@�ʑj �1-JJ�4i.�ڴR\�5�s��-v��<2��E��� 	���1MDn8<j`����n�fsn�<$F��4�����X58���\�dJ��Lr���X��]�p��zP�d�d8�w[� `�Gn��%.�F���k�[,��x���YJ]�<	�����f�y'
,��.�4��}���_!���m�+��l�3�nɻ�� Y��FD����,��*�iIZ��nY6��ـ*�>��EȐ��q��=ӿ���!Ҟg�����e���-/���@�qCs��5]O����v���/1�1�J�������f��;ᷲ�%[�Ĳ�3$a��������0R��;�*��W/B>�X���L%�3�����jA3�W�M���	�>SW�mMj\&��~L\~��va]�TE�(��,�����%�p���ix�arK���Z���**��B������Є1��/���d�@���q*�Qh+LwcA�;�:�21����  [�k�c���:u��=Fx#�{)Ө��%�&�ߧ`+��&�S���N_����jk�=$�󿆆�Xj¥:�E`�$PF�WKy1Ġ�W�X>[�$F#/��/Fw9�c�b���k1����|�@r̘�x`Ug �a洖N�q�`2�؂�^�*�G���8���!Kn�
4?'&GK��O}�҈��WUQ(�_6A?����mj=J�P8D��WJ%��lЃR�3H��C���#��!��0����i�������O1���o9	l⚒�����e��H��������P|�����CZ����L6���Ԟ�J�o]��I����U4��/����qk�Zm��*n�(����
5x!)_�D,���@h�/l�!V�A��$7ě;D~�<��C��9\Cd���>;����Řj�Vj�_+�hl���<bE,�|m$ �҉;x����K��,�H@��\q������B���r��쬚�4g�/E��	��6��eޛ�H�;���X��ߍ!��pg�L����r�4~ֈo��O�+�[��D``=�ӓ+N��=tбAe!29���S��˻s���<%�$�8e�R���76+���A�~8''��*#65�=(��u��Ʈ�A�Z�3���]>l�qd�l�+���n�'p��Cw�$�����a7'"@A;����k(2�x2�`g��%����*�m�x ��ʶ���a�R+�4Cy��<�9unqg{�_�Q3y��\�b����NN�}�Q��Ʃ�7EBʘ�:j�>�hLJq�;�p^+,ox��A��1t;�o� cy�Au��������c{�\�<MX��pG&�ش����2J8���o��`F�q�4�y�˯���yzt���?��3�S��Nl���w�/G����¢C�39dW��?�->�`?MKQ�@:h"v���U�.���]�)wf
a�vQ�K㿬�-���͖y_�F�Ƨ��t���� ��6`<���b��>]��11�; K͈]���,��L"z������+��͟��%Kboqi?��(�Ib�o�h�a!�Zy�Pѽ��v��I�t������^�M�~Y�"W`A�P�����в�+j�ɪ]-�|i�w��G�p��i�h��1���[������H��O�ަ�9ȸ���ܿ������V�i���?˩�7TچY5�r�%����߀BF�r`�ܻ\�L�]����1��T>DR�[+�hBx����%�O�!)�5C�~/�EoL��9��C�S���3�~ʿg�m;�.](�����y#�����
r3᯵Ϋ����7�����$(K��cn`W�����z��7�	.�f�W����0pʯ�[�\)	ְ'�ډ���u�>��[��C���$�Z�@���a)����O�3p���؝l�'�f}<��70Re�I��le�ԯ�F;J�ɰ? \��dE�w�&�����^k�`�s?j�Q��� _k ��۶��49�7Q$c{{{��T�b��
Gu7W��\l���y�<���n�]e�g>��k"�+���5*���qIS���s�1���a�{�,��-˪&�`���c�D�T�E�(��i:�zn��g̻A��	�1T�r4á�="d�=���V���Բ�R^����+izz߭��)�U�a���`'�YJjT�yw��(�
y7�Ս�������5���D��t�=\<:3��+([t��}�k j�D�����[�����I�v�
Cwh.�e��U��D�&VL�Rֺ� 8K;����n�_{p���)�W?��3@�*�/�[E�3�+��r9(�GK�i�#��PhF-WJg�W�5���VU�e؅aV�����n�}���E������JbC5{�YӫI��E�.�g2�ʞO'����qo,h�܁:��e��1�䌴�Ǹ��ȵ���\gS+�4��gø\��ۤ3��J�խ�)M}�i�W��o� KOg!�ޡ�楀\0���M>�o��M��ibK�I���f�5�b����~�7B䷂�#��v؞�MCp�ۥ���8a	^m����J��Z�/]��/�g~	+<�OګkE"7���'�q���qV���{��'���ȴ:���L��r�P Ȑ�a0F0ܻ�ad��d�����]'���by�O����q,�B��˂��= 1�����[�h 9ܖ�.�|�%K���s��^�f���k!� uh�>�)��W��������I�.k��}�W5��\�����7`���[�� J������L�ݾܳ�������G0�8����ֻ��^ 'Զ�u�KƦO��J�}��y�^�'[%$ڰR-B��:�-j�=���(C�,�G
�`^p}�Bt*���͏���#���ia��&��_'�F*M�ΒKϦ>�xMW_�m,#� ����jpM��0�S�am�����|�Bt-_��D��ߙ�MS7��Ol:M�0a ӡs��e����ۊ_�	�T�~wλs����U�+������%O7���'���#,Ds�����W<��j�� S	�"�T� ��7���s���v!F�n/�[o{?"�~� �	��ZF�O�%sy%ϩ0�����k皸�&�� �kG1��dP&���bC�b^/�.�ل�
�g:�\�S��$�'��Z-)�����[ F� 2�xٞ�k�%�(LʞQKTw��*�*6���2 �wu�L�
��;.Pǯ��e�;�L#�:���\bǶ�m#\ψᣗ��bp�%d/u'��͚�_�@���K�T�end�؃c�R�I�(evYY�A�#|ii���<��߿���!r�Ba����e��\�-���7�_�p����n�G���{�����XA� йI����b�v���w.[Fh���Brb_7�]?o�l�$pFn>͙g����bg�H�U$3VrNn,�B�z<[#��b��o�:O �>ǀ~��l藍���E�v�y�����e1�\W�L���u3�&'�Pa�j�V���:�A3�g�5W��<��L�ʈZ	q �L�5�d��f㛅C���Z�#S�a3z��ɲ2geb+�M�t}�t����Y2
����.�&�ۼ�V�o�>ɕN�Ǿ���V�:\��I"c
����
)�L�o��˸�2%U�?���y|��P7��Y���B�z����3��W�*�L��#�����I�� !<w�Ϡ�J��$@�R�%�ԿW��2\����t��F��i#���o�J(���b�oN��hK)}Ư�B�I�Cyxu��oP��jZ�z$T� �=��`>y���š/a�����\�;nJDɱ�bT�*[e���)+Aֻѻ�1QU�������̑�;#+�	�/X��Z�7�~���@�|�-��D��T'��yqX�{9)���o5;��ݫ������MG���<<R�x��:���i�)~�O��V&&?4P�?��BF��=�T��̞�t���Ͱp�v��M�.���(������cRA��4��c]Rm��l�E�L���^_WE�<�91b&���T8�%�H�$�:b-��3p��%�Ue�'f��R��+�(,�� ���G�G%i��F�n�,��W&�CSEh�.�u�
����1X�4�C��p����qe�Ma���-k_�Ŗ��R�.4��C�T�,�ם^����+�.$���%d[��]?ڭ�uh:�%v�ǂ�)ν�Yv&)#H�{�)�I�����nWk������)^��X���1"DVs�q2�=ˌ	��A��R����)����!':T#>��nS�����L�g��!��e�AQM�u4�	Ci�}4�|$a> (i�� ���d)7f�A7�� �>�
#�m��r� ���^�}�D���Ѡ�[�;��+B�_Z7H�$2R�,��֊�:	OF ���M��'���A�(�����WH�M�Ct'˲�ǹ�N�2$^e/�R���>M�d�qNI�%����hfB)�w>z�C%+x�BX�(�/<���1a�l	\�δ�2�Y�h�[�ʾ�Vf��z3��G<Å�Hr`���Kҥ��_ハGM�ɒK�_
�4M#~u�٤���ݵW��w��k�߮�VU+�"�2��:P9!/0�C9�?�<�N�U��}kLTD����7]�=����O�_L����?�������(����z���F`�dY�E�}	����/���U�9�x�̈́+ �$E%g�o� ��;h�ʸd&*��g��W���>�;CF��_{C���G�Y���@�称��c��c��]����Ɗ�J�#$��K�幕o:�i��?7��1*���[�3�C	i��]�ꢞ&vZ�3u����-���G6I�HND�s
_�k�T	9��J@���r�}*Y�zo�Ak��}89^�J�H�J�?���ߞo��?Bqp4{U�pF�g��o-�t����>(�e�?��y�	'0'���U�`��.���-�BN��+�f{�����t�ɬ��ϯ�a3l
�e)����nf��.T:�����zV5pIJ�L0�qi*~�8�Bn�(m�6es
q�(�B�e��a�ĳ-�&~*��M.z�0��MY/w�Z��Q���	�y���~��kb:i �ƾ��c9�Y�J�%ޞ�!���ڽr��̓���ma��ck��dz&�U�Q�^$��Y|�f�W��%�6m�P�xj��	�6m!Y`ɲ~/ q�X�,�,`�A\�l�+,NX��I�d��̓
��ٍ��kSMܢZ��E^F~��Gj2���	�'.�L�P��w�-\��t�:�� �珊�K�c[��~��m��;�'�U��]ˊ�[���oMz
���K��#sR=)̴�ѷ��6`�
(������`u8�+����U2TT��}Ơ�c-�ܚ)�^���2�*�[0^HB�Ñ屙��4w�#�DV -jjS.�E6�1T�-���R*	Iͬ�4�Pt-^���0�j�*��֜�5mR�k���"��>�Pq��lJ��w���^���5V��#�W���Ax��P=��v(�[��x��'�����u�e��"�e٠���C���c������0�|Qһ�.�>$�)9x��:ݝ����G�4$î��JS�HHt�{4cm�`���p�#G�W�4RO�tWQʰ,�؍�Y��Nt�F��WR�b��f��?���	Uw�L��E���A CI�6�;�K�2��o�[���I�_!����,$��|r�]!�6l8�@��޼8�j[]�gn�d��s�23Q�>i���b�ĉ&�ǯ��R{���J����	Y9��l���!;�ж�u}�?6� =1똅�Ob>�L)z����r��E@�|�i�A�����@A*��g��/��UX�������hydWd4 ~��juU�9��?%ZΨE�g����Q��@�����4I��ky��p5�P �AA�HKɶϖ3-��.�s�\>�e��	���;��P����s=�.襬1�l^�Ȫ������Xu�*�!�
�\�h�5��ń?�����W\A�B�4��)�T3���"x��Thpl��B��(k���e
;,�4�x8���fW��t׌ӭN�G�5��n�t�.
�By�Y���H'�.�t�e�Z�J�J�+�k9B����Ǐ���;�k�+j-��P�ZzpX.9�����s�$o���������~no+g#X�>�\���8�SΑ� ��XJ6��<p&O�4N��y��k�X����M}ѡs7m�?�2�|^�E�u���#��p�7�h�篃�nt�v����9��Ƞv>�0[����U�}.?w���ݎhp��� Ʈ�k}	u}�U2�o:";���/&5M �����i�U���6� �,��)�}ў�=��i�#�{�C~9.���_�1�Y)>qUQ�bD僱��u�?�5qZQ�B��W� }��#��{��Vp�U�ja�Q�b_U�W��X��1�:��{�1�d����V��?�ǽ�~�3:�e��� �"[�i�r��-�Fc�r�]�����.6�u�����}R�}th���a��gVIPqyb����U����^9��C~VB��w��e~C���j�.rP�{�'s�W��RG���
;�s:.8�n�5������X��|~�%��މ4����&iR�
*�V��Z��>u`,toD�NH�m8��rp���?a劮�%+ ���p�KI��ҩ�|�쪤�)�3�Ad�ȹ�S8��;v>f�4H���Gp���2���S�x�bc=���x���<oU�^�hb��������:�� �����n��
�����P�,i]t�m����O�EBE���z�5�6���l׎�������C�P�a���r�����K����t}������|�Q�������3�f���X�[�PY���[fO�?���П�"�@�8)�jӴ�r���6���˄���r6M�0�5 ��Z,���
��\��w���5r��ݴܰ�Yq���čf2��߸AA��֗|l�z��[޿�J\�(��i�*�3J/5�V?��?~��!ңy�밌��������eG�s���9إT�dDڊ��#q����D��Z�N)�s��$m�HN{?#$pd\�"x�$ʳY�~�k��s�ɝ��m�5k���Ϧ�.v݆i$��g�Q\j��!r����UT4�9<�����c�C�u��0cb�?(U�諳S����yz�49�?��*�Q؃��8E���fJc������SD"�2GC�]�Swf��V�4���p����8`ʎ6�?蘱	^���#�ek�G�2�%y��	h�K"mw �#A�ȯp�(o�ӻ��>��[��WĦ-�"��L�k�p���9J|���#�A�WW�X7�=`5�@��c�s@��c�e�V����ʘ7&ކ(�_�ܑ��'0���o����S���ӓ��,c�{����ֳ��7qd��,�i�Pq;0�g�Xʮg�l�X>�8t&��JV�5����jX��(Y�ˀS��Q4�>��H^��Yhk!�	S�kiq����u<���G��i�C�^���tg�zg%��s2}1P��S�5�[w�e�>j��lDυ˿.�����6φrω�x
Vwꚺ��DD���9��Q�aak	�gv��<!�,�_��Q_�B��y�"#rE��'^�B^a�|��{dy&�y�21n��A0���^���e֗������W`���Ni҆Ow�Ҭ�$��歎�<K�<�Z0�αJ!���h�l�K��5��'��Ѧ���v8${MVd����!����"�m�z�x���q[>��:��1�ȅ�ͅ�X���X}wR���� P��EQ����a�� gE�		%�7�(�Y{T؜�d��`�]//�W�*���~c�����1ǎ7�A~�A�[�3Iߣ�ڿ���.�<�Tn���C��
�+�����Ԭ�(?�s���4����Y�,���nW����Lr�V�}�^�FH��9S�x�
#�U���P�4O�'N����X��G<J�JP�1V�0n��QL^̲��IV�+b���6dha1�P5?����D�I�z��W���ޤ!��6B7��c�IԨ�/��_���b���X6NkG�Q!�jL��j��
��#��Ԑ�c;9:���Z ������[]/r��?����Д7oT�Aif�-C�f\/1���H�X�F�h�փ�LwP�ѝyC�s�0��d�E^�h�:�[�b�rf������s���F�jP��R7�y�XR9��^uTy�U��ZQ�0ޚ٧/�����R5zU�$ȥ��_yߴɏ�ܐ6� O'���TT�e^�Ra�V��Ķ9l�#O����oo	mw�vS��'�1<=�f�����7 �Z�T
V��GP�zA�4�>(�����P�x���񣴿�YW:��ワ�C��n�W��c��u'A��"��ih�+�ב{8��u�J���=�N���\r��ˋ����a�@���H�s�,��Kq��D���D^ᑳW�w�[*oa6����WcL��{��v�O{�����gG��V8��&	�FJ�O��2�ڤu�p<���q5�p�2� ��T<9n�LP�Ո�jIhv���Ԧ5��+� m��
8F~�)H&���\���5�=kSU!�w+Zĸ�o��$���.�WC��㏌�Q����Im2����rC���Rv�f���(\O2>cN��9+=���k�1���Zk�����q�8�<�׌���u����~�{�c�Nb�a�P�nV��Sv|̚(��l�->�(��/ը��L��vlaNʿ{���}1��3r�I�r�N���:����-o��f� ���F�H8��l��Cs�ޖ���J́�+������a�8�Ӕe�*v�#`���!��E Vn�]ܧ�C�?x�{��ꋌ�ڛys�$qi��вj)=�"M�w�%�y�����^��E��oL�<��L��߾�C���].�h�@�j��o{����Μe8PI�}<������3���!��+�
���O�EU�G��V��j���(I�[��̦�Ņie�B�%��b���2f�-d:f���= ��U1�-J�G�0ZGi��M�9��L<RW�4��OG�*��ӹ͸�A��կHl�ݏ����֐s�r�b���eg3OЫ1廏g�љĖLT��n�������PZ�h�<Q���$�Ȼ*��elL����?���������(
U����E�ѯ�c[�N�Xu��sjvs����27�R�����x_ݹp\�#����f��*�0�v�f����U�7�AL�*O.����aҗ�8��ȱ�9���3$���X�?�{x���g�{�@a���0c8�a-���+��6'J���w��2|Q�F6���[V�7��0���(j�} խ(�A{?����W�-*j41�u
%�r_�T�� �t+Wq��\�Y&��,Cq�����2ة�t��p������a���Eѥ���+2{a]��������i��*,�H-��_�q��3�xBjҥ�� 79�Q�?ś�#��c_�ڏY�i��Gx}] �t����ZY����8��}a��@=�c�"���Q����Q݋��cd��C�^�5���2(S�����K�ō��~��c��E]qE|�`��"�4�n�J�C�a�vD����_1��͜,�[�2�Z6��S��)V9��Wٞ�B��p��V6�E�DI:p��{?��k���[C�W�$�؆~a�;�n�?���֩�"�r�/p/
Ce�fE�����)�eUc>��#�ʵ���<1Ǯ�E4��N�9R'_��GF "6Z��9�V����/����O2:Y {�+�V <��h2
)�]��oĢc|�C���zߑ��d����ͼ�i�#����g.T�ɑj$3�v����nS�~)������y�*�bB�BKwvϒ̑���r�y�4E��N�����T�MS���%��8V(�ׁ�<(��~z��B����|�;�fJ�|}�s��������� ���<�N>b\����(�BT�D`B�0LDWB]���,�Ay�R:֕ＭGT�7�w$\i8G�Hc�Y������aG�8:)�[G1*�����GD!��I*�hN�}��%��M�do�	���ٓ+���ZSȅEM]���A��3E,8�B�o>8VE�� E�O����£�s"YO(]q�Ha��O���Y؁��ƍI-J�Ccy��5T	B�^��^���*� !�� e��3��S�����4=B��F�[�qR�`�q��bi8���!Y����
~�ΖT5�z����!��L(���|m��O�M> 5�cn:��� ����IF���i�('����$�R�J�H����$yf� AyG����B��00QO�+�7n�2��*N���|4˽,1��{��3]&�0l'�d	���8���5?t��
gEZ�RH���0b����z�>o�#Э��LK{1J�z�y�g�hZ����*9�-�j�s.�k=��D���-s	@���x)q ���|�Iv�~���\$�;&@����n@��RvY܃�|��2�d�БAx�yVCi�]��ѩ�pDT������ťcmԸTᬯܦ��S����{a0X~Hthm��7�l۔� �E�h�@��{9w���hZ�d[g��I? O��[�올S�������h�Bx��"7��b���x���L���Cu%Q<���$ M-g�@�͏J�X�9�u>��O��Q�����Y�7���wU�[z0�!Y�{t<o�YCc�Lc�n-�>�����[y4�F~��'�ҍgw�⌫?з�����0c�0�I����=W5j�Zػ� a[E��>г�Ɠ�;}��M͉-E����M���[c�y� �� �����ѥc9�vN�0�&�?l�_�%k�D��`��c��F���4/n�$�d�`ݑ��w�Ul�5�[�P�V�S��o�ȑH�㕷-�D���'b[Gnr@��x�mӀ���`5�1�	<��A���!�
82S��b0f���6�G4���n�~ ���؋���F�Y�.O�X���h�v6e:�,fhd)h�'$�G0o��B
�}�t��Mg�����?:��L��P��~JUUnA���"d��0�?u�O熾��6`�0�G�ú��eo����f"����3"ĆCvx:���Yҹ����� �I� ��Mh�����eCъ���.F�a�5�:�ˌ�δ=5��S�9���-%���_=,�q�33paM��l� �F�
.�ղ.q�u�?�Sc�<�np���g���j�1;\0�&X�8�2>�u���]:Y��	ܿ�e+(M�����b�{�K��;Ҵg��1]|�ݚ̓&~�՝?i�\�U���K�9��/ci
 �g&��'�@��3ق�v�Q��.6�3�N�<�|���T���(� �4�;H�9���?��ɲ��##�b(��f$�>xAx��U�ڥ7�u���fE�q����/"��BBbEߘA\�Hl�]_�֗�j��.�0;/g�x���$g��{�rU��VA3f�綃 �(��B�x�X��<���U��o��:����4�A�]\F�a_�62<r@<a��l���[-9��7�}��c�7�Ѓ@Ю�/uu���
*d
'�Μ6y&m���������ϫ�Y��<�Z_W�8#Ax�P;>J*�|����֝>����nmY���?�<�H�3vFәc���m�)G��l��^��v�
p��⏂3�
�y�\$���c��'��ww�J<IX����e9�e��^�<~BL�LQ����-J�Ɣf� �;J�O��o�ڇ���;�j�}y��a��"A֎�x�m���>�𮻇Я�[C�u����/��_����c��F����a���v�MPҽE�]w��`ˏ<�<1�Oʣ0 $yz_�G��_$��&�P����y-���D82T;�OA8E�wr��[��S+IB�Aˡ���������Y-�/bDlµ�N�5'��Ń*g��I�-g7Ǯ��ёv�D����c6�]�DO� �á�a)�q��/��舴L��p:�1�~�����@Δ��H�_��܂S����q/	I2`d_HJ�`�bݲ �T��ƛ��t��oᩯ���#�W�r�ق�*����x �f̯FX�o��<�;��/q�fl�Eo��r�֎B������1�T�X����d�4O�o���G�1X~��|(��I_:�6������SD^����I�~���B��l@��׫㩟���K���H��)����T2����!+��u�����*a�$�w�|I�!�q�39���� ��dD��9��@�����t<�/�,��`���|w���R�~�������#�� S?��40V�7Ã����.^��C��ףn+vsa%����q�iv�N{�D�P�d�7ҡa����E�g������~����Y5o�
$��]´p��.�}l3�D�F�+�50ff����'�y17ff�;�n�g+ռs�n�ɍ�L�����c���A�u$�}ٶn&��r���r^�\��%�P^�o�l�]���X����t�8���^�$[9�����:�AL۰���P��0�W��F���¿�'��{*Y��{��pxF}7@8�4T��p���&T�;C;/�B<d�z�*�R������Q�'��İ�/�Ŷ��Z:�}YS�j��o���9m�D�&;Z�ss	�n���!�!�FU��Z�����LKxI7���Xqպ��`�n�ԙ����3��-`�?��#Y�Z1迀p�^��٩m
P˔�4!��vÆՇ^
������!eLќ����i�41(\�..����?H!�NT���%M9E^�F����p�9��/�D��֮�m͠>�)r�v2�3���l��cq�L�����uSx�C���ϴ�0Ԏ���G��n��8��=�sy����X�6�iϜ�#?���Z��q�����"�y��H�/]�_k�~���Y\df����"*�tk�2�8ߙm�w	�t~c����/(+X�q{�2�C�G\�=���`L5�0^,h����'���e=
눑K���O�_��v$y�r�4��	MB�?X����g�+�����;���.f�7G�,�v$������
��4�*:N�������5����D�HaK�z�MB��	T�����C�g�v�����?'N�4Z4�L�L��(��Q}�T����(���M㝶ƈc�P(v� q�����?��1ɤ"w�]ah�O5{����7z��xˢ�H��i�va�i���~�3�Q����]�F�3_���D�2~�m^@P�ޫ�3E�}���$j�N� e�a��q� ��3T�a��Uu
`�H�!���=���x�Ǒ���{J���!�UY����?��@�,��cXPAl�e��IA��1�g^� �kQ�+z�z��������ұ��H*��J��T��j��2�4
'&	kCˇ+��P���s�=�Nޝp0.����U6��(�[�,�'��N�p̴�D<�J��
���rs�����ή�x����vUXCI5��ژ�"��mM����*�h!qE%b�/�"�K����� h��+ˣ�s�{�`��T�^	���h��Y}��K=��aoZ� ���XO���5��$T']6<�"��c�C�4Vw�c�9)|N�x��_ڼ�'/4��k󎖌f��؞�Kqps�@->Qh�L����R����8F��YֽN�뒱eݛ���~�.��T��{Q�nW<�n}�T44�� ��k 4R嫵�A�_,O�E��-gՑi/?��'(O�9�� �������y���[�2�3����s���$��N���Dq��|^��S7�|�dx��sK䫩�����8��)��kD��OX����������Uu�b�3�\�Ă�7�,tvane�Βy#)S�� �/�g�1 ����K�j�W���@a2�:��娀M����C��w�6��a�@߶}N:�t��A\l]ϖ���7�v����\q�W4AIΖ��=C�bF����ГǪn1����L˲�~�X{Fo6yn��?��"��&汄%%'����^��S�Dx�8ܥ-c
N��:<_�!�u}Z=�pG�l.݀d��!������l���i^t�j<��z�?L��T?`B2��O���X��3�ѝ���U�~k��˹�A�ݪI1V�o%�I��U��_�����@B�r�ˬ��m"O��s|r��������	�P��'�R���*���:�����Y�]��z�?Z�*6> �����U����~��d4���
nV9�ןI� ���E���]��?uH��hY����.��}�/^1K�6�8�|:��~Q�Q�K��"�8�8da��b��bpz��Q�$< ���pE��U�W
4TϜ���'�l�T�L�ۻ�����yv�-���S��<��^j͍:��z<ՊCf%DZ3>�^��v�;��O�7���	�s�U�A��!�, i�b����+���1�b)��$��G��&��(� pc���af�'�5x��^O�[�A?�31ʉ�w�ׁ�.�U��B��>���b��!C
D��@[S�Z�|�d7������eU�U=j�
�Ɍd�H,V����)��s�/�%�{l4��O��F(�?�,�\A?<�=�/\��6�&��o�_f�;dN��\a���$-Ҟ��_]E1Rh P
�� ��#yp��z�׍e/�T�Bal�������B��)-	��É�}i�nC�q,�7[����⣕��_�-�(��sՏ@�3��_��٩O��-z�^ջ�Z������L�&��A�N������'���G��$�)	e�`v���$X��$5i��<�ZE#����$��fC�~G�uZ�B�v�ä��@<i�<��?�.$[��5����?�� #��L+L�� ����ٮ�1vk[��Ir�0#Ew�A�׫Tf���-\B��el�o�� ���-��xb\��V�%ֹߵ����e�I�/����$�vfř'h�kǜW������+��oVy��OO�N��n���6I�2��,Z�l��4#�˝U΅nl�u��v<R�
;GW��E� ]X+I�o*\M��
r����`�C��Fi�������<^6�R��C=��g��c-�i����G-è2?@*���n]��G��j�LX��0^��=+�._-t�
�� 
n��\0��Ml�7#�j	�x�+���|�P!6�B=ŞA����/Ƃ{�Q�/T��9�)�UGѿ�@'Z���ٿ���#^ĕxP�[����$NƜ������'Yn �ଳ�L}���L�9�/-�v}����g��!��ӥb��� m�(h�{+� �� zxq�.]���{X%L�	W_�Y�A�.r��1�b�,F�oݤ4����RE�6R�Đ$�as����\S^���(q��~�M�r-G��3�(�	�����_j;���!ʇ����y�~w�Y4|;������*�U$����p��[���_'͋f�bw�T]a�?(�ւ��$�$�2�|�g��z�U|oZ�ۃ_�ܡ�]T�<T��{zV�a�q���Y�U���ʓ�c� ��n����!�0�s]4Uf�\�Wy����r{A�5�Q��M�0EJ5�M�n}��׏�1�/R
�t�K����"�Ӽ��"Q~5� ���5L��Eb}�@Nib�ݬ4_���,�Ơ��L	1�n7�,8@_�r껓������ͪ)ĬC��/H����?�\�QWnTF�.�]��A��a+D/ú�:w���@q��m�1}#G ~<���K:(ɒE���LP�k,��Q��;���`Z�:H����z���a�����C��.&v��bC���|����<�<OU����7}��x8$��A�Z�n�?��Rî�HY+���>|ۼBI���n\4�{{�ޅWuC���\wg���JO�Ӄ�>D�������
�h�P}�p&;!���$e�h���:�����~���L48A�g�{�/#��QRH���I�)�i��z-�TqH]
P��@�i6�Z��I�˨����^_�,�k���f񆜤� ��9��[Kl#�x �eE#ޖ��a!Cdi\�.t�7��|��� }ٯG���ݯ�`3�L5�U�Ș�'�@-�/�ٝ���Ѿ�?���qݠ�V���{���Ǚ�\�^"
�^���S��o�s����)iz�ӈO1�H��^Jf�L@�Ω���5,D��)e�C�de�NV{�/���2Ԙ:@<3v�iq䣿�f���"��{|>ޝMx�3�w�	s�TĴ��e�����F���|��F�����@"��uV���[�^���M������-
ʢ\x�U��.,�١�c�f����Ud��tb@�����
s�J��B�k���B�lV^� >.E�m��]�E�%E�%��m��{p��v��\&����R�g�Ľ3���e5�m��`~��-���K]���Z��u7[��o�ߟ}����� �{�i����h���B�}��4�1�tĲ[uh�����T��%�(�}g�@G��tΎǏ_-�ˠ)�?�`r�Т�@�3޼K�XU���JS�&�$�$U�������,�4-�%֖��|ݮ�R�<n���&�4�u�/1w�����U�jꡟ�� �,������C��̰t9�'�E�kLt4d��6 �N�ot�c���ׅ�+ܞ�bn��R|���rbtAޝx��Us�Q��v~e�ň�=��jJ2�w�X���5?=�H�"j�����qo����˻�V���Kh��>�<�A�g9�3:��JS�e�w��+�)�������CΚ��/�����Ƹ;�7���S�w�K��$��J�^ի��$��Jq�㙠�e��7� -��4�Kgj��,�I��w~$��R<��ࢅH6M��)9� ]�g����@�~�랡��sIEZ�g{-��o�wb>� ʚ������<�������'n�j��v�Oj�e�[� �L�c���r:�Q�O�Ia�55�em4���mZI!�;��d��lE��0(�����U�)�?�YQ��U����_G"%�+ak,跜l��%���0J+}H?��vD�����AV�T7*�Ϫ�!D�1���(CO��'Y�p��.����S١�R����瀟I��<�v�b�1�l}�+d��x����%�Mに�s ��=N�YB�P��\w��?+X:��)cj汐���Sx�M�'����&	S.�N	�(˱��r�Q������/n#*˧I/+,HCl�yW�j
�L�σ+�'1�!��tpl�#���B;���o\Y]PLo���7��p"��3S�D��.$
�1���	�Бp�I�r�v�N��u��e.���/���Ф+�gs�$�Z5�zv�x�U�ܖP��F��ɥk�S�W||_&O�p��,��AB|�MPvMrT�]�p�l+}ƹ[�4�Z'�}��Zw�e��Q��<��3xX ���ڊ��w�Jv&%,]|��]����Z�ll� �\�N��21E#��1���,0|;ty0
�;z��L�x��0f u
�D�/uK�Z�-*��=�z���� S��G��A���d>���������_!Eg=��H}�.� �a�(�ߞ����KR�Z�m1�wa�h��9��B�HQG���u��>${��RR#l�Z�2�a,��M��vTȇ&x��z�;3�c4o�n2$�-�P:�s#�Cj�U���(Ji��V68!�1]G� ����0��V޸[G ���)���B����R��.�$f�h�H��� ��F*9�Z�h����{H�"�ɚ ����P���$�#@�(?Y*����:R�v,�<%V�:�`LN�����$v��̘�E��:���-1{�v&�[�z���{i��F�B]��-����0G�_��=?�I�c�A�o��Ԓ�7����V�R�le����D�,b�f���	�Y�\oM�H�D�p��������Xx���%�u�~�h�LX�La�ܩ��H�:Zf0���T �J�� ��#���!&�ˆ�.*��}כ����<�!�P_E(:d������]���AJ|W��9�7;$ߡ.�
��u�e�G��	R�y�`6t\�z��O]��
�:�Itn��ߦԭ�ې�v {���|%ɈK8����g$+'���@�u|�x8%Sz��@�R�u��X��#Խ��,�'0D����W�����Ķ9e+NE�o���"��`N�A�ez�M��ҳ��'�=�]'�g�V?&0_K^G�Սb��
9�����YҙO�y� ~R��D���pO=QB�(=.O,Cndǯ�ڑ��;b�,:�������&��f�I��EM]R�O_�蠄���K����\�c�$[��|L�ITU?����\������!��$>Y�<`��y�3�l�Ai����/��vD�_ܟ���Q�4�<��	A9O�+���A��@6�@>�EY�^;��բ�����%���9�h`�x�q�hTk��[�:
f���ːc�êފ���a�-�#"2V�GM��W��L5���j�ғ�����Lx~����Ȇ�T 
^�7M�M���uF�Dw<q���h�$�3\G�!X>�Q.��"x�ǖ�
��'Iħ:tJ�1��b8�4�䧍�#qW��keLdw�M�x�l��W��]���.xv�p��~�o����� 5�K��P�
�iW�M�<&�L�\���~>ߊʖu�Us,�#u��^�Dת��x;˪0p��w7 cş��������b�>@дVj�OR�ȥ@H27 �N�$��!�x,�X�A�Ϩ}@��Ĝ6���(8o)S�IR� �N����^Pl���'m���Z8{�����_��q���f���[�̅�1��u�� ����KH`,B�� ��{�B��+��gN?���@�G��;d�k��G���/�;Qh�ړW�t�$���H%�m`<�=G�����b�癲���"��9�4x��q�y�x�P0Ap+>��o��,F�������"��p�� ���a�2��4@R�3�,�k���QN�]4i'����4cQ���32�D:~&�o��2��U����>�T�OW���OJ2/)υE��lf,V�B����G|/@h��t4���ރ����i�p�#�)t�7ю_8���V,ү&~D�-%FK��LI^��Lo��8���;'i7��{F&<Fڂ
d�)O�"�y@}��Vׯ��	_��[���c�N�ϥ{W��V��;vd���*�	�ه����Spc�$@�4��h�-�<>�s�U�[��?i�4-?_L~/��'o���ZȘ�FO���0�;���^Cʤ�xo��� <9��G��:��L�JB�z�~�9�ёZ�X�*��sQ��4w�<[�-O2���H	O��M�b���o�U.;�݇0�.1�C?��޳A��B0s"1|6�N����^ǀ{��fW}dw���AA���_��oMKɋ��b|�	�y����&��y*ɛ�"��u�%]0�y5 �C�g<#����_��>8B���!Jp;����މ�D������B-|J���H��{	}jHW��l�VZu�P�NX�m2j������/O!U�+ηcS5\F��^t>��L�&���9<���Ml}h��r��k��UK����H6XÜe������TSd��޿L�#��s�Ao���g����P�[<"g��	��P/�&�!4��+�ɕ�Y\��v��M���;i�SHβ��B~n���.�J���})��h2�ݫ+Z�v��y�$G�G�:@
=Td^U��y	�<�<�"��zf���{�[�)3��q��:�QjM�w�6�3�g�ވU��nc�7o��P�}�v�``�����I��8��mrV�i���&y9��K;�
ف`�A��e�ϭ����AO���j(����&�S�B�"�4Tf��K�	^�e<���9�r `w���=��c$VE-"�@j�/��Y.K�H�_���<�S�!���n�n�
�V���y�4�T-�b�˸�Aop���ϻ�K��6���0�~�ssu� ckQ�R�hH�2|I*��@I�!V���G�
[:A��O�,��Ԇ@N�$�|fE�_��Q���@�������Q�����:w�1\{#�۾]7(�i�'d�-����Yr����pr�'�{:p�?��މ���P��թ������>;eХX11��М�m|�C��,!L�e/"���	���>�D=^���	�@TR#��_�w��ג��rR�Uɣb������op�9ڮ�s��E��ǡ8]��A1��"8i�
�Z��kiNX�z����bI��g�]t�fM��