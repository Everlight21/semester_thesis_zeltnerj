-- DE4_QSYS.vhd

-- Generated using ACDS version 12.1sp1 243 at 2013.07.29.16:53:13

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE4_QSYS is
	port (
		spi_2_MISO                          : in    std_logic                      := '0';             --                spi_2.MISO
		spi_2_MOSI                          : out   std_logic;                                         --                     .MOSI
		spi_2_SCLK                          : out   std_logic;                                         --                     .SCLK
		spi_2_SS_n                          : out   std_logic;                                         --                     .SS_n
		spi_1_MISO                          : in    std_logic                      := '0';             --                spi_1.MISO
		spi_1_MOSI                          : out   std_logic;                                         --                     .MOSI
		spi_1_SCLK                          : out   std_logic;                                         --                     .SCLK
		spi_1_SS_n                          : out   std_logic;                                         --                     .SS_n
		dvi_master_interface_ClkDvixCI      : in    std_logic                      := '0';             -- dvi_master_interface.ClkDvixCI
		dvi_master_interface_DviNewLinexDI  : in    std_logic                      := '0';             --                     .DviNewLinexDI
		dvi_master_interface_DviNewFramexDI : in    std_logic                      := '0';             --                     .DviNewFramexDI
		dvi_master_interface_DviPixelAvxSI  : in    std_logic                      := '0';             --                     .DviPixelAvxSI
		dvi_master_interface_DviDataOutxDO  : out   std_logic_vector(31 downto 0);                     --                     .DviDataOutxDO
		oct_rdn                             : in    std_logic                      := '0';             --                  oct.rdn
		oct_rup                             : in    std_logic                      := '0';             --                     .rup
		no_of_cam_channels_export           : out   std_logic_vector(3 downto 0);                      --   no_of_cam_channels.export
		led_export                          : out   std_logic_vector(7 downto 0);                      --                  led.export
		button_export                       : in    std_logic_vector(3 downto 0)   := (others => '0'); --               button.export
		reset_reset_n                       : in    std_logic                      := '0';             --                reset.reset_n
		clk_clk                             : in    std_logic                      := '0';             --                  clk.clk
		cmv_master_interface_PixelValidxSI  : in    std_logic                      := '0';             -- cmv_master_interface.PixelValidxSI
		cmv_master_interface_RowValidxSI    : in    std_logic                      := '0';             --                     .RowValidxSI
		cmv_master_interface_FrameValidxSI  : in    std_logic                      := '0';             --                     .FrameValidxSI
		cmv_master_interface_DataInxDI      : in    std_logic_vector(159 downto 0) := (others => '0'); --                     .DataInxDI
		cmv_master_interface_ClkLvdsRxxCI   : in    std_logic                      := '0';             --                     .ClkLvdsRxxCI
		memory_mem_a                        : out   std_logic_vector(13 downto 0);                     --               memory.mem_a
		memory_mem_ba                       : out   std_logic_vector(2 downto 0);                      --                     .mem_ba
		memory_mem_ck                       : out   std_logic_vector(1 downto 0);                      --                     .mem_ck
		memory_mem_ck_n                     : out   std_logic_vector(1 downto 0);                      --                     .mem_ck_n
		memory_mem_cke                      : out   std_logic_vector(0 downto 0);                      --                     .mem_cke
		memory_mem_cs_n                     : out   std_logic_vector(0 downto 0);                      --                     .mem_cs_n
		memory_mem_dm                       : out   std_logic_vector(7 downto 0);                      --                     .mem_dm
		memory_mem_ras_n                    : out   std_logic_vector(0 downto 0);                      --                     .mem_ras_n
		memory_mem_cas_n                    : out   std_logic_vector(0 downto 0);                      --                     .mem_cas_n
		memory_mem_we_n                     : out   std_logic_vector(0 downto 0);                      --                     .mem_we_n
		memory_mem_dq                       : inout std_logic_vector(63 downto 0)  := (others => '0'); --                     .mem_dq
		memory_mem_dqs                      : inout std_logic_vector(7 downto 0)   := (others => '0'); --                     .mem_dqs
		memory_mem_dqs_n                    : inout std_logic_vector(7 downto 0)   := (others => '0'); --                     .mem_dqs_n
		memory_mem_odt                      : out   std_logic_vector(0 downto 0)                       --                     .mem_odt
	);
end entity DE4_QSYS;

architecture rtl of DE4_QSYS is
	component DE4_QSYS_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			clken      : in  std_logic                     := 'X';             -- clken
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X'              -- reset
		);
	end component DE4_QSYS_onchip_memory;

	component DE4_QSYS_mem_if_ddr2_emif is
		port (
			pll_ref_clk       : in    std_logic                      := 'X';             -- clk
			global_reset_n    : in    std_logic                      := 'X';             -- reset_n
			soft_reset_n      : in    std_logic                      := 'X';             -- reset_n
			afi_clk           : out   std_logic;                                         -- clk
			afi_half_clk      : out   std_logic;                                         -- clk
			afi_reset_n       : out   std_logic;                                         -- reset_n
			mem_a             : out   std_logic_vector(13 downto 0);                     -- mem_a
			mem_ba            : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck            : out   std_logic_vector(1 downto 0);                      -- mem_ck
			mem_ck_n          : out   std_logic_vector(1 downto 0);                      -- mem_ck_n
			mem_cke           : out   std_logic_vector(0 downto 0);                      -- mem_cke
			mem_cs_n          : out   std_logic_vector(0 downto 0);                      -- mem_cs_n
			mem_dm            : out   std_logic_vector(7 downto 0);                      -- mem_dm
			mem_ras_n         : out   std_logic_vector(0 downto 0);                      -- mem_ras_n
			mem_cas_n         : out   std_logic_vector(0 downto 0);                      -- mem_cas_n
			mem_we_n          : out   std_logic_vector(0 downto 0);                      -- mem_we_n
			mem_dq            : inout std_logic_vector(63 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs           : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n         : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt           : out   std_logic_vector(0 downto 0);                      -- mem_odt
			avl_ready         : out   std_logic;                                         -- waitrequest_n
			avl_burstbegin    : in    std_logic                      := 'X';             -- beginbursttransfer
			avl_addr          : in    std_logic_vector(24 downto 0)  := (others => 'X'); -- address
			avl_rdata_valid   : out   std_logic;                                         -- readdatavalid
			avl_rdata         : out   std_logic_vector(255 downto 0);                    -- readdata
			avl_wdata         : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avl_be            : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req      : in    std_logic                      := 'X';             -- read
			avl_write_req     : in    std_logic                      := 'X';             -- write
			avl_size          : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			local_init_done   : out   std_logic;                                         -- local_init_done
			local_cal_success : out   std_logic;                                         -- local_cal_success
			local_cal_fail    : out   std_logic;                                         -- local_cal_fail
			oct_rdn           : in    std_logic                      := 'X';             -- rdn
			oct_rup           : in    std_logic                      := 'X'              -- rup
		);
	end component DE4_QSYS_mem_if_ddr2_emif;

	component DE4_QSYS_nios2_qsys is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(30 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                          : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(18 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_begintransfer       : in  std_logic                     := 'X';             -- begintransfer
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_select              : in  std_logic                     := 'X';             -- chipselect
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component DE4_QSYS_nios2_qsys;

	component DE4_QSYS_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DE4_QSYS_jtag_uart;

	component DE4_QSYS_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DE4_QSYS_sysid;

	component DE4_QSYS_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DE4_QSYS_timer;

	component DE4_QSYS_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component DE4_QSYS_led;

	component DE4_QSYS_button is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component DE4_QSYS_button;

	component DE4_QSYS_mm_clock_crossing_bridge_io is
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(9 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component DE4_QSYS_mm_clock_crossing_bridge_io;

	component DE4_QSYS_spi_2 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component DE4_QSYS_spi_2;

	component DE4_QSYS_no_of_cam_channels is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component DE4_QSYS_no_of_cam_channels;

	component DE4_QSYS_cmv_master_interface_0 is
		port (
			ClkxCI          : in  std_logic                      := 'X';             -- clk
			RstxRBI         : in  std_logic                      := 'X';             -- reset_n
			AMWritexSO      : out std_logic;                                         -- write
			AMWriteDataxDO  : out std_logic_vector(127 downto 0);                    -- writedata
			AMAddressxDO    : out std_logic_vector(31 downto 0);                     -- address
			AMBurstCountxSO : out std_logic_vector(7 downto 0);                      -- burstcount
			AMWaitReqxSI    : in  std_logic                      := 'X';             -- waitrequest
			PixelValidxSI   : in  std_logic                      := 'X';             -- export
			RowValidxSI     : in  std_logic                      := 'X';             -- export
			FrameValidxSI   : in  std_logic                      := 'X';             -- export
			DataInxDI       : in  std_logic_vector(159 downto 0) := (others => 'X'); -- export
			ClkLvdsRxxCI    : in  std_logic                      := 'X'              -- export
		);
	end component DE4_QSYS_cmv_master_interface_0;

	component DE4_QSYS_dvi_master_interface_0 is
		port (
			ClkxCI             : in  std_logic                     := 'X';             -- clk
			RstxRBI            : in  std_logic                     := 'X';             -- reset_n
			AmWaitReqxSI       : in  std_logic                     := 'X';             -- waitrequest
			AmAddressxDO       : out std_logic_vector(31 downto 0);                    -- address
			AmReadDataxDI      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			AmReadxSO          : out std_logic;                                        -- read
			AmReadDataValidxSI : in  std_logic                     := 'X';             -- readdatavalid
			AmBurstCountxDO    : out std_logic_vector(7 downto 0);                     -- burstcount
			ClkDvixCI          : in  std_logic                     := 'X';             -- export
			DviNewLinexDI      : in  std_logic                     := 'X';             -- export
			DviNewFramexDI     : in  std_logic                     := 'X';             -- export
			DviPixelAvxSI      : in  std_logic                     := 'X';             -- export
			DviDataOutxDO      : out std_logic_vector(31 downto 0)                     -- export
		);
	end component DE4_QSYS_dvi_master_interface_0;

	component DE4_QSYS_nios2_qsys_instruction_master_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid  : out std_logic                                         -- readdatavalid
		);
	end component DE4_QSYS_nios2_qsys_instruction_master_translator;

	component DE4_QSYS_nios2_qsys_data_master_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(5 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_burstcount     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid  : out std_logic;                                        -- readdatavalid
			av_write          : in  std_logic                     := 'X';             -- write
			av_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess    : in  std_logic                     := 'X'              -- debugaccess
		);
	end component DE4_QSYS_nios2_qsys_data_master_translator;

	component DE4_QSYS_mm_clock_crossing_bridge_io_m0_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_burstcount     : in  std_logic                     := 'X';             -- burstcount
			av_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid  : out std_logic;                                        -- readdatavalid
			av_write          : in  std_logic                     := 'X';             -- write
			av_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess    : in  std_logic                     := 'X'              -- debugaccess
		);
	end component DE4_QSYS_mm_clock_crossing_bridge_io_m0_translator;

	component DE4_QSYS_dvi_master_interface_0_avalon_master_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(9 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_burstcount     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid  : out std_logic                                         -- readdatavalid
		);
	end component DE4_QSYS_dvi_master_interface_0_avalon_master_translator;

	component DE4_QSYS_cmv_master_interface_0_avalon_master_translator is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			uav_address       : out std_logic_vector(31 downto 0);                     -- address
			uav_burstcount    : out std_logic_vector(11 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                         -- read
			uav_write         : out std_logic;                                         -- write
			uav_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(15 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(127 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                         -- lock
			uav_debugaccess   : out std_logic;                                         -- debugaccess
			av_address        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                         -- waitrequest
			av_burstcount     : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			av_write          : in  std_logic                      := 'X';             -- write
			av_writedata      : in  std_logic_vector(127 downto 0) := (others => 'X')  -- writedata
		);
	end component DE4_QSYS_cmv_master_interface_0_avalon_master_translator;

	component DE4_QSYS_nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			av_address       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write         : in  std_logic                      := 'X';             -- write
			av_read          : in  std_logic                      := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest   : out std_logic;                                         -- waitrequest
			av_readdatavalid : out std_logic;                                         -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                      := 'X';             -- debugaccess
			av_lock          : in  std_logic                      := 'X';             -- lock
			cp_valid         : out std_logic;                                         -- valid
			cp_data          : out std_logic_vector(126 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                         -- startofpacket
			cp_endofpacket   : out std_logic;                                         -- endofpacket
			cp_ready         : in  std_logic                      := 'X';             -- ready
			rp_valid         : in  std_logic                      := 'X';             -- valid
			rp_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rp_ready         : out std_logic                                          -- ready
		);
	end component DE4_QSYS_nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent;

	component DE4_QSYS_nios2_qsys_data_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			av_address       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write         : in  std_logic                      := 'X';             -- write
			av_read          : in  std_logic                      := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest   : out std_logic;                                         -- waitrequest
			av_readdatavalid : out std_logic;                                         -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                      := 'X';             -- debugaccess
			av_lock          : in  std_logic                      := 'X';             -- lock
			cp_valid         : out std_logic;                                         -- valid
			cp_data          : out std_logic_vector(126 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                         -- startofpacket
			cp_endofpacket   : out std_logic;                                         -- endofpacket
			cp_ready         : in  std_logic                      := 'X';             -- ready
			rp_valid         : in  std_logic                      := 'X';             -- valid
			rp_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rp_ready         : out std_logic                                          -- ready
		);
	end component DE4_QSYS_nios2_qsys_data_master_translator_avalon_universal_master_0_agent;

	component DE4_QSYS_mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			av_address       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write         : in  std_logic                      := 'X';             -- write
			av_read          : in  std_logic                      := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest   : out std_logic;                                         -- waitrequest
			av_readdatavalid : out std_logic;                                         -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                      := 'X';             -- debugaccess
			av_lock          : in  std_logic                      := 'X';             -- lock
			cp_valid         : out std_logic;                                         -- valid
			cp_data          : out std_logic_vector(126 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                         -- startofpacket
			cp_endofpacket   : out std_logic;                                         -- endofpacket
			cp_ready         : in  std_logic                      := 'X';             -- ready
			rp_valid         : in  std_logic                      := 'X';             -- valid
			rp_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rp_ready         : out std_logic                                          -- ready
		);
	end component DE4_QSYS_mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent;

	component DE4_QSYS_dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			av_address       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write         : in  std_logic                      := 'X';             -- write
			av_read          : in  std_logic                      := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest   : out std_logic;                                         -- waitrequest
			av_readdatavalid : out std_logic;                                         -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                      := 'X';             -- debugaccess
			av_lock          : in  std_logic                      := 'X';             -- lock
			cp_valid         : out std_logic;                                         -- valid
			cp_data          : out std_logic_vector(126 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                         -- startofpacket
			cp_endofpacket   : out std_logic;                                         -- endofpacket
			cp_ready         : in  std_logic                      := 'X';             -- ready
			rp_valid         : in  std_logic                      := 'X';             -- valid
			rp_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rp_ready         : out std_logic                                          -- ready
		);
	end component DE4_QSYS_dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent;

	component DE4_QSYS_cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			av_address       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write         : in  std_logic                      := 'X';             -- write
			av_read          : in  std_logic                      := 'X';             -- read
			av_writedata     : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(127 downto 0);                    -- readdata
			av_waitrequest   : out std_logic;                                         -- waitrequest
			av_readdatavalid : out std_logic;                                         -- readdatavalid
			av_byteenable    : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                      := 'X';             -- debugaccess
			av_lock          : in  std_logic                      := 'X';             -- lock
			cp_valid         : out std_logic;                                         -- valid
			cp_data          : out std_logic_vector(234 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                         -- startofpacket
			cp_endofpacket   : out std_logic;                                         -- endofpacket
			cp_ready         : in  std_logic                      := 'X';             -- ready
			rp_valid         : in  std_logic                      := 'X';             -- valid
			rp_data          : in  std_logic_vector(234 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rp_ready         : out std_logic                                          -- ready
		);
	end component DE4_QSYS_cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent;

	component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(127 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component DE4_QSYS_onchip_memory_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_onchip_memory_s1_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(127 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			in_data   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid  : in  std_logic                     := 'X';             -- valid
			in_ready  : out std_logic;                                        -- ready
			out_data  : out std_logic_vector(31 downto 0);                    -- data
			out_valid : out std_logic;                                        -- valid
			out_ready : in  std_logic                     := 'X'              -- ready
		);
	end component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			in_data   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid  : in  std_logic                     := 'X';             -- valid
			in_ready  : out std_logic;                                        -- ready
			out_data  : out std_logic_vector(31 downto 0);                    -- data
			out_valid : out std_logic;                                        -- valid
			out_ready : in  std_logic                     := 'X'              -- ready
		);
	end component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component DE4_QSYS_led_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_led_s1_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_timer_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_timer_s1_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_spi_2_spi_control_port_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_spi_2_spi_control_port_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_sysid_control_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_sysid_control_slave_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(12 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(255 downto 0);                    -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(378 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(379 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(379 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(255 downto 0)                     -- data
		);
	end component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(379 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(379 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo is
		port (
			clk       : in  std_logic                      := 'X';             -- clk
			reset     : in  std_logic                      := 'X';             -- reset
			in_data   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			in_valid  : in  std_logic                      := 'X';             -- valid
			in_ready  : out std_logic;                                         -- ready
			out_data  : out std_logic_vector(255 downto 0);                    -- data
			out_valid : out std_logic;                                         -- valid
			out_ready : in  std_logic                      := 'X'              -- ready
		);
	end component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component DE4_QSYS_spi_1_spi_control_port_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_spi_1_spi_control_port_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(126 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(127 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component DE4_QSYS_no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent;

	component DE4_QSYS_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(126 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_addr_router;

	component DE4_QSYS_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(126 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_addr_router_001;

	component DE4_QSYS_addr_router_002 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(126 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_addr_router_002;

	component DE4_QSYS_addr_router_003 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(126 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_addr_router_003;

	component DE4_QSYS_addr_router_004 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(234 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(234 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_addr_router_004;

	component DE4_QSYS_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(126 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_id_router;

	component DE4_QSYS_id_router_002 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(126 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_id_router_002;

	component DE4_QSYS_id_router_004 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(126 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_id_router_004;

	component DE4_QSYS_id_router_009 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(378 downto 0);                    -- data
			src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_id_router_009;

	component DE4_QSYS_limiter is
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(126 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(126 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(11 downto 0)                      -- data
		);
	end component DE4_QSYS_limiter;

	component DE4_QSYS_limiter_001 is
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(126 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(126 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(11 downto 0)                      -- data
		);
	end component DE4_QSYS_limiter_001;

	component DE4_QSYS_limiter_002 is
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(126 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(126 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(11 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(11 downto 0)                      -- data
		);
	end component DE4_QSYS_limiter_002;

	component DE4_QSYS_burst_adapter is
		port (
			clk                   : in  std_logic                      := 'X';             -- clk
			reset                 : in  std_logic                      := 'X';             -- reset
			sink0_valid           : in  std_logic                      := 'X';             -- valid
			sink0_data            : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                         -- ready
			source0_valid         : out std_logic;                                         -- valid
			source0_data          : out std_logic_vector(126 downto 0);                    -- data
			source0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			source0_startofpacket : out std_logic;                                         -- startofpacket
			source0_endofpacket   : out std_logic;                                         -- endofpacket
			source0_ready         : in  std_logic                      := 'X'              -- ready
		);
	end component DE4_QSYS_burst_adapter;

	component DE4_QSYS_burst_adapter_002 is
		port (
			clk                   : in  std_logic                      := 'X';             -- clk
			reset                 : in  std_logic                      := 'X';             -- reset
			sink0_valid           : in  std_logic                      := 'X';             -- valid
			sink0_data            : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                         -- ready
			source0_valid         : out std_logic;                                         -- valid
			source0_data          : out std_logic_vector(126 downto 0);                    -- data
			source0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			source0_startofpacket : out std_logic;                                         -- startofpacket
			source0_endofpacket   : out std_logic;                                         -- endofpacket
			source0_ready         : in  std_logic                      := 'X'              -- ready
		);
	end component DE4_QSYS_burst_adapter_002;

	component DE4_QSYS_rst_controller is
		port (
			reset_in0 : in  std_logic := 'X'; -- reset
			clk       : in  std_logic := 'X'; -- clk
			reset_out : out std_logic         -- reset
		);
	end component DE4_QSYS_rst_controller;

	component DE4_QSYS_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(126 downto 0);                    -- data
			src0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(126 downto 0);                    -- data
			src1_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_cmd_xbar_demux;

	component DE4_QSYS_cmd_xbar_demux_001 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			sink_ready          : out std_logic;                                         -- ready
			sink_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- data
			src0_ready          : in  std_logic                      := 'X';             -- ready
			src0_valid          : out std_logic;                                         -- valid
			src0_data           : out std_logic_vector(126 downto 0);                    -- data
			src0_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src0_startofpacket  : out std_logic;                                         -- startofpacket
			src0_endofpacket    : out std_logic;                                         -- endofpacket
			src1_ready          : in  std_logic                      := 'X';             -- ready
			src1_valid          : out std_logic;                                         -- valid
			src1_data           : out std_logic_vector(126 downto 0);                    -- data
			src1_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src1_startofpacket  : out std_logic;                                         -- startofpacket
			src1_endofpacket    : out std_logic;                                         -- endofpacket
			src2_ready          : in  std_logic                      := 'X';             -- ready
			src2_valid          : out std_logic;                                         -- valid
			src2_data           : out std_logic_vector(126 downto 0);                    -- data
			src2_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src2_startofpacket  : out std_logic;                                         -- startofpacket
			src2_endofpacket    : out std_logic;                                         -- endofpacket
			src3_ready          : in  std_logic                      := 'X';             -- ready
			src3_valid          : out std_logic;                                         -- valid
			src3_data           : out std_logic_vector(126 downto 0);                    -- data
			src3_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src3_startofpacket  : out std_logic;                                         -- startofpacket
			src3_endofpacket    : out std_logic;                                         -- endofpacket
			src4_ready          : in  std_logic                      := 'X';             -- ready
			src4_valid          : out std_logic;                                         -- valid
			src4_data           : out std_logic_vector(126 downto 0);                    -- data
			src4_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src4_startofpacket  : out std_logic;                                         -- startofpacket
			src4_endofpacket    : out std_logic;                                         -- endofpacket
			src5_ready          : in  std_logic                      := 'X';             -- ready
			src5_valid          : out std_logic;                                         -- valid
			src5_data           : out std_logic_vector(126 downto 0);                    -- data
			src5_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src5_startofpacket  : out std_logic;                                         -- startofpacket
			src5_endofpacket    : out std_logic;                                         -- endofpacket
			src6_ready          : in  std_logic                      := 'X';             -- ready
			src6_valid          : out std_logic;                                         -- valid
			src6_data           : out std_logic_vector(126 downto 0);                    -- data
			src6_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src6_startofpacket  : out std_logic;                                         -- startofpacket
			src6_endofpacket    : out std_logic;                                         -- endofpacket
			src7_ready          : in  std_logic                      := 'X';             -- ready
			src7_valid          : out std_logic;                                         -- valid
			src7_data           : out std_logic_vector(126 downto 0);                    -- data
			src7_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src7_startofpacket  : out std_logic;                                         -- startofpacket
			src7_endofpacket    : out std_logic;                                         -- endofpacket
			src8_ready          : in  std_logic                      := 'X';             -- ready
			src8_valid          : out std_logic;                                         -- valid
			src8_data           : out std_logic_vector(126 downto 0);                    -- data
			src8_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src8_startofpacket  : out std_logic;                                         -- startofpacket
			src8_endofpacket    : out std_logic;                                         -- endofpacket
			src9_ready          : in  std_logic                      := 'X';             -- ready
			src9_valid          : out std_logic;                                         -- valid
			src9_data           : out std_logic_vector(126 downto 0);                    -- data
			src9_channel        : out std_logic_vector(11 downto 0);                     -- channel
			src9_startofpacket  : out std_logic;                                         -- startofpacket
			src9_endofpacket    : out std_logic;                                         -- endofpacket
			src10_ready         : in  std_logic                      := 'X';             -- ready
			src10_valid         : out std_logic;                                         -- valid
			src10_data          : out std_logic_vector(126 downto 0);                    -- data
			src10_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src10_startofpacket : out std_logic;                                         -- startofpacket
			src10_endofpacket   : out std_logic;                                         -- endofpacket
			src11_ready         : in  std_logic                      := 'X';             -- ready
			src11_valid         : out std_logic;                                         -- valid
			src11_data          : out std_logic_vector(126 downto 0);                    -- data
			src11_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src11_startofpacket : out std_logic;                                         -- startofpacket
			src11_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_cmd_xbar_demux_001;

	component DE4_QSYS_cmd_xbar_demux_002 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(126 downto 0);                    -- data
			src0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(126 downto 0);                    -- data
			src1_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(126 downto 0);                    -- data
			src2_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic;                                         -- endofpacket
			src3_ready         : in  std_logic                      := 'X';             -- ready
			src3_valid         : out std_logic;                                         -- valid
			src3_data          : out std_logic_vector(126 downto 0);                    -- data
			src3_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                         -- startofpacket
			src3_endofpacket   : out std_logic;                                         -- endofpacket
			src4_ready         : in  std_logic                      := 'X';             -- ready
			src4_valid         : out std_logic;                                         -- valid
			src4_data          : out std_logic_vector(126 downto 0);                    -- data
			src4_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                         -- startofpacket
			src4_endofpacket   : out std_logic;                                         -- endofpacket
			src5_ready         : in  std_logic                      := 'X';             -- ready
			src5_valid         : out std_logic;                                         -- valid
			src5_data          : out std_logic_vector(126 downto 0);                    -- data
			src5_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src5_startofpacket : out std_logic;                                         -- startofpacket
			src5_endofpacket   : out std_logic;                                         -- endofpacket
			src6_ready         : in  std_logic                      := 'X';             -- ready
			src6_valid         : out std_logic;                                         -- valid
			src6_data          : out std_logic_vector(126 downto 0);                    -- data
			src6_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src6_startofpacket : out std_logic;                                         -- startofpacket
			src6_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_cmd_xbar_demux_002;

	component DE4_QSYS_cmd_xbar_demux_003 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(126 downto 0);                    -- data
			src0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_cmd_xbar_demux_003;

	component DE4_QSYS_cmd_xbar_demux_004 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(234 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(234 downto 0);                    -- data
			src0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_cmd_xbar_demux_004;

	component DE4_QSYS_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(126 downto 0);                    -- data
			src_channel         : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component DE4_QSYS_cmd_xbar_mux;

	component DE4_QSYS_cmd_xbar_mux_009 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(378 downto 0);                    -- data
			src_channel         : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component DE4_QSYS_cmd_xbar_mux_009;

	component DE4_QSYS_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(126 downto 0);                    -- data
			src0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(126 downto 0);                    -- data
			src1_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_rsp_xbar_demux;

	component DE4_QSYS_rsp_xbar_demux_009 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(378 downto 0);                    -- data
			src0_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(378 downto 0);                    -- data
			src1_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(378 downto 0);                    -- data
			src2_channel       : out std_logic_vector(11 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component DE4_QSYS_rsp_xbar_demux_009;

	component DE4_QSYS_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(126 downto 0);                    -- data
			src_channel         : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component DE4_QSYS_rsp_xbar_mux;

	component DE4_QSYS_rsp_xbar_mux_001 is
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			src_ready            : in  std_logic                      := 'X';             -- ready
			src_valid            : out std_logic;                                         -- valid
			src_data             : out std_logic_vector(126 downto 0);                    -- data
			src_channel          : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket    : out std_logic;                                         -- startofpacket
			src_endofpacket      : out std_logic;                                         -- endofpacket
			sink0_ready          : out std_logic;                                         -- ready
			sink0_valid          : in  std_logic                      := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                         -- ready
			sink1_valid          : in  std_logic                      := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                         -- ready
			sink2_valid          : in  std_logic                      := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                         -- ready
			sink3_valid          : in  std_logic                      := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                         -- ready
			sink4_valid          : in  std_logic                      := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                         -- ready
			sink5_valid          : in  std_logic                      := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                         -- ready
			sink6_valid          : in  std_logic                      := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                         -- ready
			sink7_valid          : in  std_logic                      := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                         -- ready
			sink8_valid          : in  std_logic                      := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                         -- ready
			sink9_valid          : in  std_logic                      := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                         -- ready
			sink10_valid         : in  std_logic                      := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                         -- ready
			sink11_valid         : in  std_logic                      := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component DE4_QSYS_rsp_xbar_mux_001;

	component DE4_QSYS_rsp_xbar_mux_002 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(126 downto 0);                    -- data
			src_channel         : out std_logic_vector(11 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                         -- ready
			sink3_valid         : in  std_logic                      := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                         -- ready
			sink4_valid         : in  std_logic                      := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                         -- ready
			sink5_valid         : in  std_logic                      := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                         -- ready
			sink6_valid         : in  std_logic                      := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component DE4_QSYS_rsp_xbar_mux_002;

	component DE4_QSYS_width_adapter is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_ready          : out std_logic;                                         -- ready
			in_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_data          : out std_logic_vector(378 downto 0);                    -- data
			out_channel       : out std_logic_vector(11 downto 0);                     -- channel
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic                                          -- startofpacket
		);
	end component DE4_QSYS_width_adapter;

	component DE4_QSYS_width_adapter_002 is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_ready          : out std_logic;                                         -- ready
			in_data           : in  std_logic_vector(234 downto 0) := (others => 'X'); -- data
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_data          : out std_logic_vector(378 downto 0);                    -- data
			out_channel       : out std_logic_vector(11 downto 0);                     -- channel
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic                                          -- startofpacket
		);
	end component DE4_QSYS_width_adapter_002;

	component DE4_QSYS_width_adapter_003 is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_ready          : out std_logic;                                         -- ready
			in_data           : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_data          : out std_logic_vector(126 downto 0);                    -- data
			out_channel       : out std_logic_vector(11 downto 0);                     -- channel
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic                                          -- startofpacket
		);
	end component DE4_QSYS_width_adapter_003;

	component DE4_QSYS_width_adapter_005 is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_ready          : out std_logic;                                         -- ready
			in_data           : in  std_logic_vector(378 downto 0) := (others => 'X'); -- data
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_data          : out std_logic_vector(234 downto 0);                    -- data
			out_channel       : out std_logic_vector(11 downto 0);                     -- channel
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic                                          -- startofpacket
		);
	end component DE4_QSYS_width_adapter_005;

	component DE4_QSYS_crosser is
		port (
			in_clk            : in  std_logic                      := 'X';             -- clk
			in_reset          : in  std_logic                      := 'X';             -- reset
			out_clk           : in  std_logic                      := 'X';             -- clk
			out_reset         : in  std_logic                      := 'X';             -- reset
			in_ready          : out std_logic;                                         -- ready
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_channel        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- channel
			in_data           : in  std_logic_vector(126 downto 0) := (others => 'X'); -- data
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_valid         : out std_logic;                                         -- valid
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_channel       : out std_logic_vector(11 downto 0);                     -- channel
			out_data          : out std_logic_vector(126 downto 0)                     -- data
		);
	end component DE4_QSYS_crosser;

	component DE4_QSYS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DE4_QSYS_irq_mapper;

	component DE4_QSYS_irq_synchronizer is
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component DE4_QSYS_irq_synchronizer;

	component de4_qsys_nios2_qsys_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(8 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect         : out std_logic;                                        -- chipselect
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_read               : out std_logic;                                        -- read
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component de4_qsys_nios2_qsys_jtag_debug_module_translator;

	component de4_qsys_onchip_memory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(14 downto 0);                    -- address
			av_write              : out std_logic;                                        -- write
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			av_read               : out std_logic;                                        -- read
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component de4_qsys_onchip_memory_s1_translator;

	component de4_qsys_jtag_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(0 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect         : out std_logic;                                        -- chipselect
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable    : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component de4_qsys_jtag_uart_avalon_jtag_slave_translator;

	component de4_qsys_mm_clock_crossing_bridge_io_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(9 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component de4_qsys_mm_clock_crossing_bridge_io_s0_translator;

	component de4_qsys_button_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(1 downto 0);                     -- address
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component de4_qsys_button_s1_translator;

	component de4_qsys_timer_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(2 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_readdata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect         : out std_logic;                                        -- chipselect
			av_read               : out std_logic;                                        -- read
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component de4_qsys_timer_s1_translator;

	component de4_qsys_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(0 downto 0);                     -- address
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component de4_qsys_sysid_control_slave_translator;

	component de4_qsys_mem_if_ddr2_emif_avl_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                      := 'X';             -- clk
			reset                 : in  std_logic                      := 'X';             -- reset
			uav_address           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(12 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                      := 'X';             -- read
			uav_write             : in  std_logic                      := 'X';             -- write
			uav_waitrequest       : out std_logic;                                         -- waitrequest
			uav_readdatavalid     : out std_logic;                                         -- readdatavalid
			uav_byteenable        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(255 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                      := 'X';             -- lock
			uav_debugaccess       : in  std_logic                      := 'X';             -- debugaccess
			av_address            : out std_logic_vector(24 downto 0);                     -- address
			av_write              : out std_logic;                                         -- write
			av_read               : out std_logic;                                         -- read
			av_readdata           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(255 downto 0);                    -- writedata
			av_beginbursttransfer : out std_logic;                                         -- beginbursttransfer
			av_burstcount         : out std_logic_vector(7 downto 0);                      -- burstcount
			av_byteenable         : out std_logic_vector(31 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                      := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			av_begintransfer      : out std_logic;                                         -- begintransfer
			av_writebyteenable    : out std_logic_vector(31 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                         -- lock
			av_chipselect         : out std_logic;                                         -- chipselect
			av_clken              : out std_logic;                                         -- clken
			uav_clken             : in  std_logic                      := 'X';             -- clken
			av_debugaccess        : out std_logic;                                         -- debugaccess
			av_outputenable       : out std_logic                                          -- outputenable
		);
	end component de4_qsys_mem_if_ddr2_emif_avl_translator;

	signal mem_if_ddr2_emif_afi_clk_clk                                                                        : std_logic;                      -- mem_if_ddr2_emif:afi_clk -> [addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_009:clk, cmv_master_interface_0:ClkxCI, cmv_master_interface_0_avalon_master_translator:clk, cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:clk, crosser:in_clk, crosser_001:in_clk, crosser_002:in_clk, crosser_003:in_clk, crosser_004:in_clk, crosser_005:in_clk, crosser_006:in_clk, crosser_007:in_clk, crosser_008:in_clk, crosser_009:in_clk, crosser_010:in_clk, crosser_011:in_clk, crosser_012:in_clk, crosser_013:in_clk, crosser_014:in_clk, crosser_015:out_clk, crosser_016:out_clk, crosser_017:out_clk, crosser_018:out_clk, crosser_019:out_clk, crosser_020:out_clk, crosser_021:out_clk, crosser_022:out_clk, crosser_023:out_clk, crosser_024:out_clk, crosser_025:out_clk, crosser_026:out_clk, crosser_027:out_clk, crosser_028:out_clk, crosser_029:out_clk, dvi_master_interface_0:ClkxCI, dvi_master_interface_0_avalon_master_translator:clk, dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_009:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, limiter_002:clk, mem_if_ddr2_emif_avl_translator:clk, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:clk, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, mm_clock_crossing_bridge_io:m0_clk, mm_clock_crossing_bridge_io_m0_translator:clk, mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:clk, nios2_qsys:clk, nios2_qsys_data_master_translator:clk, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_instruction_master_translator:clk, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_jtag_debug_module_translator:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory:clk, onchip_memory_s1_translator:clk, onchip_memory_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_009:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_002:clk, rst_controller:clk, rst_controller_002:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk]
	signal nios2_qsys_instruction_master_waitrequest                                                           : std_logic;                      -- nios2_qsys_instruction_master_translator:av_waitrequest -> nios2_qsys:i_waitrequest
	signal nios2_qsys_instruction_master_address                                                               : std_logic_vector(18 downto 0);  -- nios2_qsys:i_address -> nios2_qsys_instruction_master_translator:av_address
	signal nios2_qsys_instruction_master_read                                                                  : std_logic;                      -- nios2_qsys:i_read -> nios2_qsys_instruction_master_translator:av_read
	signal nios2_qsys_instruction_master_readdata                                                              : std_logic_vector(31 downto 0);  -- nios2_qsys_instruction_master_translator:av_readdata -> nios2_qsys:i_readdata
	signal nios2_qsys_instruction_master_readdatavalid                                                         : std_logic;                      -- nios2_qsys_instruction_master_translator:av_readdatavalid -> nios2_qsys:i_readdatavalid
	signal nios2_qsys_data_master_burstcount                                                                   : std_logic_vector(3 downto 0);   -- nios2_qsys:d_burstcount -> nios2_qsys_data_master_translator:av_burstcount
	signal nios2_qsys_data_master_waitrequest                                                                  : std_logic;                      -- nios2_qsys_data_master_translator:av_waitrequest -> nios2_qsys:d_waitrequest
	signal nios2_qsys_data_master_writedata                                                                    : std_logic_vector(31 downto 0);  -- nios2_qsys:d_writedata -> nios2_qsys_data_master_translator:av_writedata
	signal nios2_qsys_data_master_address                                                                      : std_logic_vector(30 downto 0);  -- nios2_qsys:d_address -> nios2_qsys_data_master_translator:av_address
	signal nios2_qsys_data_master_write                                                                        : std_logic;                      -- nios2_qsys:d_write -> nios2_qsys_data_master_translator:av_write
	signal nios2_qsys_data_master_read                                                                         : std_logic;                      -- nios2_qsys:d_read -> nios2_qsys_data_master_translator:av_read
	signal nios2_qsys_data_master_readdata                                                                     : std_logic_vector(31 downto 0);  -- nios2_qsys_data_master_translator:av_readdata -> nios2_qsys:d_readdata
	signal nios2_qsys_data_master_debugaccess                                                                  : std_logic;                      -- nios2_qsys:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_data_master_translator:av_debugaccess
	signal nios2_qsys_data_master_readdatavalid                                                                : std_logic;                      -- nios2_qsys_data_master_translator:av_readdatavalid -> nios2_qsys:d_readdatavalid
	signal nios2_qsys_data_master_byteenable                                                                   : std_logic_vector(3 downto 0);   -- nios2_qsys:d_byteenable -> nios2_qsys_data_master_translator:av_byteenable
	signal mm_clock_crossing_bridge_io_m0_burstcount                                                           : std_logic_vector(0 downto 0);   -- mm_clock_crossing_bridge_io:m0_burstcount -> mm_clock_crossing_bridge_io_m0_translator:av_burstcount
	signal mm_clock_crossing_bridge_io_m0_waitrequest                                                          : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator:av_waitrequest -> mm_clock_crossing_bridge_io:m0_waitrequest
	signal mm_clock_crossing_bridge_io_m0_address                                                              : std_logic_vector(9 downto 0);   -- mm_clock_crossing_bridge_io:m0_address -> mm_clock_crossing_bridge_io_m0_translator:av_address
	signal mm_clock_crossing_bridge_io_m0_writedata                                                            : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io:m0_writedata -> mm_clock_crossing_bridge_io_m0_translator:av_writedata
	signal mm_clock_crossing_bridge_io_m0_write                                                                : std_logic;                      -- mm_clock_crossing_bridge_io:m0_write -> mm_clock_crossing_bridge_io_m0_translator:av_write
	signal mm_clock_crossing_bridge_io_m0_read                                                                 : std_logic;                      -- mm_clock_crossing_bridge_io:m0_read -> mm_clock_crossing_bridge_io_m0_translator:av_read
	signal mm_clock_crossing_bridge_io_m0_readdata                                                             : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_m0_translator:av_readdata -> mm_clock_crossing_bridge_io:m0_readdata
	signal mm_clock_crossing_bridge_io_m0_debugaccess                                                          : std_logic;                      -- mm_clock_crossing_bridge_io:m0_debugaccess -> mm_clock_crossing_bridge_io_m0_translator:av_debugaccess
	signal mm_clock_crossing_bridge_io_m0_byteenable                                                           : std_logic_vector(3 downto 0);   -- mm_clock_crossing_bridge_io:m0_byteenable -> mm_clock_crossing_bridge_io_m0_translator:av_byteenable
	signal mm_clock_crossing_bridge_io_m0_readdatavalid                                                        : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator:av_readdatavalid -> mm_clock_crossing_bridge_io:m0_readdatavalid
	signal dvi_master_interface_0_avalon_master_burstcount                                                     : std_logic_vector(7 downto 0);   -- dvi_master_interface_0:AmBurstCountxDO -> dvi_master_interface_0_avalon_master_translator:av_burstcount
	signal dvi_master_interface_0_avalon_master_waitrequest                                                    : std_logic;                      -- dvi_master_interface_0_avalon_master_translator:av_waitrequest -> dvi_master_interface_0:AmWaitReqxSI
	signal dvi_master_interface_0_avalon_master_address                                                        : std_logic_vector(31 downto 0);  -- dvi_master_interface_0:AmAddressxDO -> dvi_master_interface_0_avalon_master_translator:av_address
	signal dvi_master_interface_0_avalon_master_read                                                           : std_logic;                      -- dvi_master_interface_0:AmReadxSO -> dvi_master_interface_0_avalon_master_translator:av_read
	signal dvi_master_interface_0_avalon_master_readdata                                                       : std_logic_vector(31 downto 0);  -- dvi_master_interface_0_avalon_master_translator:av_readdata -> dvi_master_interface_0:AmReadDataxDI
	signal dvi_master_interface_0_avalon_master_readdatavalid                                                  : std_logic;                      -- dvi_master_interface_0_avalon_master_translator:av_readdatavalid -> dvi_master_interface_0:AmReadDataValidxSI
	signal cmv_master_interface_0_avalon_master_waitrequest                                                    : std_logic;                      -- cmv_master_interface_0_avalon_master_translator:av_waitrequest -> cmv_master_interface_0:AMWaitReqxSI
	signal cmv_master_interface_0_avalon_master_burstcount                                                     : std_logic_vector(7 downto 0);   -- cmv_master_interface_0:AMBurstCountxSO -> cmv_master_interface_0_avalon_master_translator:av_burstcount
	signal cmv_master_interface_0_avalon_master_address                                                        : std_logic_vector(31 downto 0);  -- cmv_master_interface_0:AMAddressxDO -> cmv_master_interface_0_avalon_master_translator:av_address
	signal cmv_master_interface_0_avalon_master_writedata                                                      : std_logic_vector(127 downto 0); -- cmv_master_interface_0:AMWriteDataxDO -> cmv_master_interface_0_avalon_master_translator:av_writedata
	signal cmv_master_interface_0_avalon_master_write                                                          : std_logic;                      -- cmv_master_interface_0:AMWritexSO -> cmv_master_interface_0_avalon_master_translator:av_write
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata                               : std_logic_vector(31 downto 0);  -- nios2_qsys_jtag_debug_module_translator:av_writedata -> nios2_qsys:jtag_debug_module_writedata
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address                                 : std_logic_vector(8 downto 0);   -- nios2_qsys_jtag_debug_module_translator:av_address -> nios2_qsys:jtag_debug_module_address
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect                              : std_logic;                      -- nios2_qsys_jtag_debug_module_translator:av_chipselect -> nios2_qsys:jtag_debug_module_select
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write                                   : std_logic;                      -- nios2_qsys_jtag_debug_module_translator:av_write -> nios2_qsys:jtag_debug_module_write
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                : std_logic_vector(31 downto 0);  -- nios2_qsys:jtag_debug_module_readdata -> nios2_qsys_jtag_debug_module_translator:av_readdata
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer                           : std_logic;                      -- nios2_qsys_jtag_debug_module_translator:av_begintransfer -> nios2_qsys:jtag_debug_module_begintransfer
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                             : std_logic;                      -- nios2_qsys_jtag_debug_module_translator:av_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                              : std_logic_vector(3 downto 0);   -- nios2_qsys_jtag_debug_module_translator:av_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	signal onchip_memory_s1_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator:av_writedata -> onchip_memory:writedata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_address                                             : std_logic_vector(14 downto 0);  -- onchip_memory_s1_translator:av_address -> onchip_memory:address
	signal onchip_memory_s1_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                      -- onchip_memory_s1_translator:av_chipselect -> onchip_memory:chipselect
	signal onchip_memory_s1_translator_avalon_anti_slave_0_clken                                               : std_logic;                      -- onchip_memory_s1_translator:av_clken -> onchip_memory:clken
	signal onchip_memory_s1_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- onchip_memory_s1_translator:av_write -> onchip_memory:write
	signal onchip_memory_s1_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(31 downto 0);  -- onchip_memory:readdata -> onchip_memory_s1_translator:av_readdata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_byteenable                                          : std_logic_vector(3 downto 0);   -- onchip_memory_s1_translator:av_byteenable -> onchip_memory:byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                              : std_logic;                      -- jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                  : std_logic_vector(0 downto 0);   -- jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                      -- mm_clock_crossing_bridge_io:s0_waitrequest -> mm_clock_crossing_bridge_io_s0_translator:av_waitrequest
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_burstcount                            : std_logic_vector(0 downto 0);   -- mm_clock_crossing_bridge_io_s0_translator:av_burstcount -> mm_clock_crossing_bridge_io:s0_burstcount
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_s0_translator:av_writedata -> mm_clock_crossing_bridge_io:s0_writedata
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_address                               : std_logic_vector(9 downto 0);   -- mm_clock_crossing_bridge_io_s0_translator:av_address -> mm_clock_crossing_bridge_io:s0_address
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator:av_write -> mm_clock_crossing_bridge_io:s0_write
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator:av_read -> mm_clock_crossing_bridge_io:s0_read
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io:s0_readdata -> mm_clock_crossing_bridge_io_s0_translator:av_readdata
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator:av_debugaccess -> mm_clock_crossing_bridge_io:s0_debugaccess
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdatavalid                         : std_logic;                      -- mm_clock_crossing_bridge_io:s0_readdatavalid -> mm_clock_crossing_bridge_io_s0_translator:av_readdatavalid
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- mm_clock_crossing_bridge_io_s0_translator:av_byteenable -> mm_clock_crossing_bridge_io:s0_byteenable
	signal button_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);   -- button_s1_translator:av_address -> button:address
	signal button_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0);  -- button:readdata -> button_s1_translator:av_readdata
	signal led_s1_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(31 downto 0);  -- led_s1_translator:av_writedata -> led:writedata
	signal led_s1_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(1 downto 0);   -- led_s1_translator:av_address -> led:address
	signal led_s1_translator_avalon_anti_slave_0_chipselect                                                    : std_logic;                      -- led_s1_translator:av_chipselect -> led:chipselect
	signal led_s1_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- led_s1_translator:av_write -> led_s1_translator_avalon_anti_slave_0_write:in
	signal led_s1_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(31 downto 0);  -- led:readdata -> led_s1_translator:av_readdata
	signal timer_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(15 downto 0);  -- timer_s1_translator:av_writedata -> timer:writedata
	signal timer_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(2 downto 0);   -- timer_s1_translator:av_address -> timer:address
	signal timer_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                      -- timer_s1_translator:av_chipselect -> timer:chipselect
	signal timer_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- timer_s1_translator:av_write -> timer_s1_translator_avalon_anti_slave_0_write:in
	signal timer_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(15 downto 0);  -- timer:readdata -> timer_s1_translator:av_readdata
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_writedata                                     : std_logic_vector(15 downto 0);  -- spi_2_spi_control_port_translator:av_writedata -> spi_2:data_from_cpu
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_address                                       : std_logic_vector(2 downto 0);   -- spi_2_spi_control_port_translator:av_address -> spi_2:mem_addr
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_chipselect                                    : std_logic;                      -- spi_2_spi_control_port_translator:av_chipselect -> spi_2:spi_select
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_write                                         : std_logic;                      -- spi_2_spi_control_port_translator:av_write -> spi_2_spi_control_port_translator_avalon_anti_slave_0_write:in
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_read                                          : std_logic;                      -- spi_2_spi_control_port_translator:av_read -> spi_2_spi_control_port_translator_avalon_anti_slave_0_read:in
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_readdata                                      : std_logic_vector(15 downto 0);  -- spi_2:data_to_cpu -> spi_2_spi_control_port_translator:av_readdata
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                          : std_logic_vector(0 downto 0);   -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(31 downto 0);  -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal mem_if_ddr2_emif_avl_waitrequest                                                                    : std_logic;                      -- mem_if_ddr2_emif:avl_ready -> mem_if_ddr2_emif_avl_waitrequest:in
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_burstcount                                      : std_logic_vector(7 downto 0);   -- mem_if_ddr2_emif_avl_translator:av_burstcount -> mem_if_ddr2_emif:avl_size
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_writedata                                       : std_logic_vector(255 downto 0); -- mem_if_ddr2_emif_avl_translator:av_writedata -> mem_if_ddr2_emif:avl_wdata
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_address                                         : std_logic_vector(24 downto 0);  -- mem_if_ddr2_emif_avl_translator:av_address -> mem_if_ddr2_emif:avl_addr
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_write                                           : std_logic;                      -- mem_if_ddr2_emif_avl_translator:av_write -> mem_if_ddr2_emif:avl_write_req
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_beginbursttransfer                              : std_logic;                      -- mem_if_ddr2_emif_avl_translator:av_beginbursttransfer -> mem_if_ddr2_emif:avl_burstbegin
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_read                                            : std_logic;                      -- mem_if_ddr2_emif_avl_translator:av_read -> mem_if_ddr2_emif:avl_read_req
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdata                                        : std_logic_vector(255 downto 0); -- mem_if_ddr2_emif:avl_rdata -> mem_if_ddr2_emif_avl_translator:av_readdata
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdatavalid                                   : std_logic;                      -- mem_if_ddr2_emif:avl_rdata_valid -> mem_if_ddr2_emif_avl_translator:av_readdatavalid
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_byteenable                                      : std_logic_vector(31 downto 0);  -- mem_if_ddr2_emif_avl_translator:av_byteenable -> mem_if_ddr2_emif:avl_be
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_writedata                                     : std_logic_vector(15 downto 0);  -- spi_1_spi_control_port_translator:av_writedata -> spi_1:data_from_cpu
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_address                                       : std_logic_vector(2 downto 0);   -- spi_1_spi_control_port_translator:av_address -> spi_1:mem_addr
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_chipselect                                    : std_logic;                      -- spi_1_spi_control_port_translator:av_chipselect -> spi_1:spi_select
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_write                                         : std_logic;                      -- spi_1_spi_control_port_translator:av_write -> spi_1_spi_control_port_translator_avalon_anti_slave_0_write:in
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_read                                          : std_logic;                      -- spi_1_spi_control_port_translator:av_read -> spi_1_spi_control_port_translator_avalon_anti_slave_0_read:in
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_readdata                                      : std_logic_vector(15 downto 0);  -- spi_1:data_to_cpu -> spi_1_spi_control_port_translator:av_readdata
	signal no_of_cam_channels_s1_translator_avalon_anti_slave_0_writedata                                      : std_logic_vector(31 downto 0);  -- no_of_cam_channels_s1_translator:av_writedata -> no_of_cam_channels:writedata
	signal no_of_cam_channels_s1_translator_avalon_anti_slave_0_address                                        : std_logic_vector(1 downto 0);   -- no_of_cam_channels_s1_translator:av_address -> no_of_cam_channels:address
	signal no_of_cam_channels_s1_translator_avalon_anti_slave_0_chipselect                                     : std_logic;                      -- no_of_cam_channels_s1_translator:av_chipselect -> no_of_cam_channels:chipselect
	signal no_of_cam_channels_s1_translator_avalon_anti_slave_0_write                                          : std_logic;                      -- no_of_cam_channels_s1_translator:av_write -> no_of_cam_channels_s1_translator_avalon_anti_slave_0_write:in
	signal no_of_cam_channels_s1_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0);  -- no_of_cam_channels:readdata -> no_of_cam_channels_s1_translator:av_readdata
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest                      : std_logic;                      -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_instruction_master_translator:uav_waitrequest
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount                       : std_logic_vector(2 downto 0);   -- nios2_qsys_instruction_master_translator:uav_burstcount -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata                        : std_logic_vector(31 downto 0);  -- nios2_qsys_instruction_master_translator:uav_writedata -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_address                          : std_logic_vector(31 downto 0);  -- nios2_qsys_instruction_master_translator:uav_address -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock                             : std_logic;                      -- nios2_qsys_instruction_master_translator:uav_lock -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_write                            : std_logic;                      -- nios2_qsys_instruction_master_translator:uav_write -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_read                             : std_logic;                      -- nios2_qsys_instruction_master_translator:uav_read -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata                         : std_logic_vector(31 downto 0);  -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_instruction_master_translator:uav_readdata
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess                      : std_logic;                      -- nios2_qsys_instruction_master_translator:uav_debugaccess -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable                       : std_logic_vector(3 downto 0);   -- nios2_qsys_instruction_master_translator:uav_byteenable -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid                    : std_logic;                      -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_instruction_master_translator:uav_readdatavalid
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest                             : std_logic;                      -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_data_master_translator:uav_waitrequest
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount                              : std_logic_vector(5 downto 0);   -- nios2_qsys_data_master_translator:uav_burstcount -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_writedata                               : std_logic_vector(31 downto 0);  -- nios2_qsys_data_master_translator:uav_writedata -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_address                                 : std_logic_vector(31 downto 0);  -- nios2_qsys_data_master_translator:uav_address -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_lock                                    : std_logic;                      -- nios2_qsys_data_master_translator:uav_lock -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_write                                   : std_logic;                      -- nios2_qsys_data_master_translator:uav_write -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_read                                    : std_logic;                      -- nios2_qsys_data_master_translator:uav_read -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_readdata                                : std_logic_vector(31 downto 0);  -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_data_master_translator:uav_readdata
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess                             : std_logic;                      -- nios2_qsys_data_master_translator:uav_debugaccess -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable                              : std_logic_vector(3 downto 0);   -- nios2_qsys_data_master_translator:uav_byteenable -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid                           : std_logic;                      -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_data_master_translator:uav_readdatavalid
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_waitrequest                     : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> mm_clock_crossing_bridge_io_m0_translator:uav_waitrequest
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_burstcount                      : std_logic_vector(2 downto 0);   -- mm_clock_crossing_bridge_io_m0_translator:uav_burstcount -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_burstcount
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_writedata                       : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_m0_translator:uav_writedata -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_writedata
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_address                         : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_m0_translator:uav_address -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_address
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_lock                            : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator:uav_lock -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_lock
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_write                           : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator:uav_write -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_write
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_read                            : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator:uav_read -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_read
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdata                        : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_readdata -> mm_clock_crossing_bridge_io_m0_translator:uav_readdata
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_debugaccess                     : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator:uav_debugaccess -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_byteenable                      : std_logic_vector(3 downto 0);   -- mm_clock_crossing_bridge_io_m0_translator:uav_byteenable -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_byteenable
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdatavalid                   : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> mm_clock_crossing_bridge_io_m0_translator:uav_readdatavalid
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_waitrequest               : std_logic;                      -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dvi_master_interface_0_avalon_master_translator:uav_waitrequest
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_burstcount                : std_logic_vector(9 downto 0);   -- dvi_master_interface_0_avalon_master_translator:uav_burstcount -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_writedata                 : std_logic_vector(31 downto 0);  -- dvi_master_interface_0_avalon_master_translator:uav_writedata -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_address                   : std_logic_vector(31 downto 0);  -- dvi_master_interface_0_avalon_master_translator:uav_address -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_lock                      : std_logic;                      -- dvi_master_interface_0_avalon_master_translator:uav_lock -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_write                     : std_logic;                      -- dvi_master_interface_0_avalon_master_translator:uav_write -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_read                      : std_logic;                      -- dvi_master_interface_0_avalon_master_translator:uav_read -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdata                  : std_logic_vector(31 downto 0);  -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> dvi_master_interface_0_avalon_master_translator:uav_readdata
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_debugaccess               : std_logic;                      -- dvi_master_interface_0_avalon_master_translator:uav_debugaccess -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_byteenable                : std_logic_vector(3 downto 0);   -- dvi_master_interface_0_avalon_master_translator:uav_byteenable -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid             : std_logic;                      -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dvi_master_interface_0_avalon_master_translator:uav_readdatavalid
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_waitrequest               : std_logic;                      -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cmv_master_interface_0_avalon_master_translator:uav_waitrequest
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_burstcount                : std_logic_vector(11 downto 0);  -- cmv_master_interface_0_avalon_master_translator:uav_burstcount -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_writedata                 : std_logic_vector(127 downto 0); -- cmv_master_interface_0_avalon_master_translator:uav_writedata -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_address                   : std_logic_vector(31 downto 0);  -- cmv_master_interface_0_avalon_master_translator:uav_address -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_lock                      : std_logic;                      -- cmv_master_interface_0_avalon_master_translator:uav_lock -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_write                     : std_logic;                      -- cmv_master_interface_0_avalon_master_translator:uav_write -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_read                      : std_logic;                      -- cmv_master_interface_0_avalon_master_translator:uav_read -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdata                  : std_logic_vector(127 downto 0); -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> cmv_master_interface_0_avalon_master_translator:uav_readdata
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_debugaccess               : std_logic;                      -- cmv_master_interface_0_avalon_master_translator:uav_debugaccess -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_byteenable                : std_logic_vector(15 downto 0);  -- cmv_master_interface_0_avalon_master_translator:uav_byteenable -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid             : std_logic;                      -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cmv_master_interface_0_avalon_master_translator:uav_readdatavalid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest               : std_logic;                      -- nios2_qsys_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                : std_logic_vector(2 downto 0);   -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_jtag_debug_module_translator:uav_burstcount
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                 : std_logic_vector(31 downto 0);  -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_jtag_debug_module_translator:uav_writedata
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                   : std_logic_vector(31 downto 0);  -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_jtag_debug_module_translator:uav_address
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                     : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_jtag_debug_module_translator:uav_write
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                      : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_jtag_debug_module_translator:uav_lock
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                      : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_jtag_debug_module_translator:uav_read
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                  : std_logic_vector(31 downto 0);  -- nios2_qsys_jtag_debug_module_translator:uav_readdata -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid             : std_logic;                      -- nios2_qsys_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess               : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_jtag_debug_module_translator:uav_debugaccess
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                : std_logic_vector(3 downto 0);   -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_jtag_debug_module_translator:uav_byteenable
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket        : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid              : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket      : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data               : std_logic_vector(127 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready              : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket     : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid           : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket   : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data            : std_logic_vector(127 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready           : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid         : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data          : std_logic_vector(31 downto 0);  -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready         : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                           : std_logic;                      -- onchip_memory_s1_translator:uav_waitrequest -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                            : std_logic_vector(2 downto 0);   -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_s1_translator:uav_burstcount
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata                             : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_s1_translator:uav_writedata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address                               : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_s1_translator:uav_address
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write                                 : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_s1_translator:uav_write
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock                                  : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_s1_translator:uav_lock
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read                                  : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_s1_translator:uav_read
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata                              : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator:uav_readdata -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                         : std_logic;                      -- onchip_memory_s1_translator:uav_readdatavalid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                           : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_s1_translator:uav_debugaccess
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                            : std_logic_vector(3 downto 0);   -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_s1_translator:uav_byteenable
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                    : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                          : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                  : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data                           : std_logic_vector(127 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                          : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                 : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                       : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket               : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                        : std_logic_vector(127 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                       : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                     : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                      : std_logic_vector(31 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                     : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(127 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(127 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator:uav_waitrequest -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> mm_clock_crossing_bridge_io_s0_translator:uav_burstcount
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> mm_clock_crossing_bridge_io_s0_translator:uav_writedata
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_address -> mm_clock_crossing_bridge_io_s0_translator:uav_address
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_write -> mm_clock_crossing_bridge_io_s0_translator:uav_write
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_lock -> mm_clock_crossing_bridge_io_s0_translator:uav_lock
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_read -> mm_clock_crossing_bridge_io_s0_translator:uav_read
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_s0_translator:uav_readdata -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator:uav_readdatavalid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mm_clock_crossing_bridge_io_s0_translator:uav_debugaccess
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> mm_clock_crossing_bridge_io_s0_translator:uav_byteenable
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(127 downto 0); -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(127 downto 0); -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid       : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data        : std_logic_vector(31 downto 0);  -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready       : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                      -- button_s1_translator:uav_waitrequest -> button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);   -- button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_s1_translator:uav_burstcount
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0);  -- button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_s1_translator:uav_writedata
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(31 downto 0);  -- button_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_s1_translator:uav_address
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_s1_translator:uav_write
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_s1_translator:uav_lock
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_s1_translator:uav_read
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0);  -- button_s1_translator:uav_readdata -> button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                      -- button_s1_translator:uav_readdatavalid -> button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_s1_translator:uav_debugaccess
	signal button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);   -- button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_s1_translator:uav_byteenable
	signal button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal button_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(127 downto 0); -- button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(127 downto 0); -- button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(31 downto 0);  -- button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                            : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                             : std_logic_vector(31 downto 0);  -- button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                            : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(2 downto 0);   -- led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(31 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(31 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(31 downto 0);  -- led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(3 downto 0);   -- led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(127 downto 0); -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(127 downto 0); -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(31 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                               : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                : std_logic_vector(31 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                               : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(31 downto 0);  -- timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(127 downto 0); -- timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(127 downto 0); -- timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(31 downto 0);  -- timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                             : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                              : std_logic_vector(31 downto 0);  -- timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                             : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest                     : std_logic;                      -- spi_2_spi_control_port_translator:uav_waitrequest -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount                      : std_logic_vector(2 downto 0);   -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> spi_2_spi_control_port_translator:uav_burstcount
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata                       : std_logic_vector(31 downto 0);  -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> spi_2_spi_control_port_translator:uav_writedata
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address                         : std_logic_vector(31 downto 0);  -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> spi_2_spi_control_port_translator:uav_address
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write                           : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> spi_2_spi_control_port_translator:uav_write
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock                            : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> spi_2_spi_control_port_translator:uav_lock
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read                            : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> spi_2_spi_control_port_translator:uav_read
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata                        : std_logic_vector(31 downto 0);  -- spi_2_spi_control_port_translator:uav_readdata -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid                   : std_logic;                      -- spi_2_spi_control_port_translator:uav_readdatavalid -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess                     : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spi_2_spi_control_port_translator:uav_debugaccess
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable                      : std_logic_vector(3 downto 0);   -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> spi_2_spi_control_port_translator:uav_byteenable
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket              : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid                    : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket            : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data                     : std_logic_vector(127 downto 0); -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready                    : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket           : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                 : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket         : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                  : std_logic_vector(127 downto 0); -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                 : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid               : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                : std_logic_vector(31 downto 0);  -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready               : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid               : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                : std_logic_vector(31 downto 0);  -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready               : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(127 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(127 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                   : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest                       : std_logic;                      -- mem_if_ddr2_emif_avl_translator:uav_waitrequest -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_burstcount                        : std_logic_vector(12 downto 0);  -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> mem_if_ddr2_emif_avl_translator:uav_burstcount
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_writedata                         : std_logic_vector(255 downto 0); -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> mem_if_ddr2_emif_avl_translator:uav_writedata
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_address                           : std_logic_vector(31 downto 0);  -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_address -> mem_if_ddr2_emif_avl_translator:uav_address
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_write                             : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_write -> mem_if_ddr2_emif_avl_translator:uav_write
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_lock                              : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_lock -> mem_if_ddr2_emif_avl_translator:uav_lock
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_read                              : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_read -> mem_if_ddr2_emif_avl_translator:uav_read
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdata                          : std_logic_vector(255 downto 0); -- mem_if_ddr2_emif_avl_translator:uav_readdata -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid                     : std_logic;                      -- mem_if_ddr2_emif_avl_translator:uav_readdatavalid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess                       : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mem_if_ddr2_emif_avl_translator:uav_debugaccess
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_byteenable                        : std_logic_vector(31 downto 0);  -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> mem_if_ddr2_emif_avl_translator:uav_byteenable
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_valid                      : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket              : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_data                       : std_logic_vector(379 downto 0); -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_ready                      : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket             : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                   : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket           : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                    : std_logic_vector(379 downto 0); -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                   : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                 : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                  : std_logic_vector(255 downto 0); -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                 : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                 : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                  : std_logic_vector(255 downto 0); -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                 : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest                     : std_logic;                      -- spi_1_spi_control_port_translator:uav_waitrequest -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount                      : std_logic_vector(2 downto 0);   -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> spi_1_spi_control_port_translator:uav_burstcount
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata                       : std_logic_vector(31 downto 0);  -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> spi_1_spi_control_port_translator:uav_writedata
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address                         : std_logic_vector(31 downto 0);  -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> spi_1_spi_control_port_translator:uav_address
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write                           : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> spi_1_spi_control_port_translator:uav_write
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock                            : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> spi_1_spi_control_port_translator:uav_lock
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read                            : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> spi_1_spi_control_port_translator:uav_read
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata                        : std_logic_vector(31 downto 0);  -- spi_1_spi_control_port_translator:uav_readdata -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid                   : std_logic;                      -- spi_1_spi_control_port_translator:uav_readdatavalid -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess                     : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spi_1_spi_control_port_translator:uav_debugaccess
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable                      : std_logic_vector(3 downto 0);   -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> spi_1_spi_control_port_translator:uav_byteenable
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket              : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid                    : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket            : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data                     : std_logic_vector(127 downto 0); -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready                    : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket           : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                 : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket         : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                  : std_logic_vector(127 downto 0); -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                 : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid               : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                : std_logic_vector(31 downto 0);  -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready               : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid               : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                : std_logic_vector(31 downto 0);  -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready               : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                      -- no_of_cam_channels_s1_translator:uav_waitrequest -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);   -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> no_of_cam_channels_s1_translator:uav_burstcount
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0);  -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> no_of_cam_channels_s1_translator:uav_writedata
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(31 downto 0);  -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_address -> no_of_cam_channels_s1_translator:uav_address
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_write -> no_of_cam_channels_s1_translator:uav_write
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_lock -> no_of_cam_channels_s1_translator:uav_lock
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_read -> no_of_cam_channels_s1_translator:uav_read
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0);  -- no_of_cam_channels_s1_translator:uav_readdata -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                      -- no_of_cam_channels_s1_translator:uav_readdatavalid -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> no_of_cam_channels_s1_translator:uav_debugaccess
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);   -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> no_of_cam_channels_s1_translator:uav_byteenable
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(127 downto 0); -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(127 downto 0); -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(31 downto 0);  -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                 : std_logic_vector(31 downto 0);  -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket             : std_logic;                      -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                   : std_logic;                      -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket           : std_logic;                      -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data                    : std_logic_vector(126 downto 0); -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                   : std_logic;                      -- addr_router:sink_ready -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                    : std_logic;                      -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid                          : std_logic;                      -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                  : std_logic;                      -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data                           : std_logic_vector(126 downto 0); -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready                          : std_logic;                      -- addr_router_001:sink_ready -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket            : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_valid                  : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket          : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_data                   : std_logic_vector(126 downto 0); -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	signal mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_ready                  : std_logic;                      -- addr_router_002:sink_ready -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_ready
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket      : std_logic;                      -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid            : std_logic;                      -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket    : std_logic;                      -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data             : std_logic_vector(126 downto 0); -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	signal dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready            : std_logic;                      -- addr_router_003:sink_ready -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket      : std_logic;                      -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid            : std_logic;                      -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket    : std_logic;                      -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data             : std_logic_vector(234 downto 0); -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	signal cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready            : std_logic;                      -- addr_router_004:sink_ready -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket               : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                     : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket             : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                      : std_logic_vector(126 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                     : std_logic;                      -- id_router:sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                           : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid                                 : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                         : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data                                  : std_logic_vector(126 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready                                 : std_logic;                      -- id_router_001:sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(126 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(126 downto 0); -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_003:sink_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal button_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal button_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(126 downto 0); -- button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal button_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                      -- id_router_004:sink_ready -> button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(126 downto 0); -- led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_005:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(126 downto 0); -- timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_006:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket                     : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid                           : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket                   : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data                            : std_logic_vector(126 downto 0); -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready                           : std_logic;                      -- id_router_007:sink_ready -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(126 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_008:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket                       : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_valid                             : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket                     : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_data                              : std_logic_vector(378 downto 0); -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_ready                             : std_logic;                      -- id_router_009:sink_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_ready
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket                     : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid                           : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket                   : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data                            : std_logic_vector(126 downto 0); -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready                           : std_logic;                      -- id_router_010:sink_ready -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(126 downto 0); -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                      -- id_router_011:sink_ready -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                         : std_logic;                      -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                               : std_logic;                      -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                       : std_logic;                      -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                                : std_logic_vector(126 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                             : std_logic_vector(11 downto 0);  -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                               : std_logic;                      -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                         : std_logic;                      -- limiter:rsp_src_endofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                               : std_logic;                      -- limiter:rsp_src_valid -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                       : std_logic;                      -- limiter:rsp_src_startofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                                : std_logic_vector(126 downto 0); -- limiter:rsp_src_data -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                             : std_logic_vector(11 downto 0);  -- limiter:rsp_src_channel -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                               : std_logic;                      -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal addr_router_001_src_endofpacket                                                                     : std_logic;                      -- addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	signal addr_router_001_src_valid                                                                           : std_logic;                      -- addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	signal addr_router_001_src_startofpacket                                                                   : std_logic;                      -- addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	signal addr_router_001_src_data                                                                            : std_logic_vector(126 downto 0); -- addr_router_001:src_data -> limiter_001:cmd_sink_data
	signal addr_router_001_src_channel                                                                         : std_logic_vector(11 downto 0);  -- addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	signal addr_router_001_src_ready                                                                           : std_logic;                      -- limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	signal limiter_001_rsp_src_endofpacket                                                                     : std_logic;                      -- limiter_001:rsp_src_endofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_001_rsp_src_valid                                                                           : std_logic;                      -- limiter_001:rsp_src_valid -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_001_rsp_src_startofpacket                                                                   : std_logic;                      -- limiter_001:rsp_src_startofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_001_rsp_src_data                                                                            : std_logic_vector(126 downto 0); -- limiter_001:rsp_src_data -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_001_rsp_src_channel                                                                         : std_logic_vector(11 downto 0);  -- limiter_001:rsp_src_channel -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_001_rsp_src_ready                                                                           : std_logic;                      -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	signal addr_router_002_src_endofpacket                                                                     : std_logic;                      -- addr_router_002:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	signal addr_router_002_src_valid                                                                           : std_logic;                      -- addr_router_002:src_valid -> limiter_002:cmd_sink_valid
	signal addr_router_002_src_startofpacket                                                                   : std_logic;                      -- addr_router_002:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	signal addr_router_002_src_data                                                                            : std_logic_vector(126 downto 0); -- addr_router_002:src_data -> limiter_002:cmd_sink_data
	signal addr_router_002_src_channel                                                                         : std_logic_vector(11 downto 0);  -- addr_router_002:src_channel -> limiter_002:cmd_sink_channel
	signal addr_router_002_src_ready                                                                           : std_logic;                      -- limiter_002:cmd_sink_ready -> addr_router_002:src_ready
	signal limiter_002_rsp_src_endofpacket                                                                     : std_logic;                      -- limiter_002:rsp_src_endofpacket -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_002_rsp_src_valid                                                                           : std_logic;                      -- limiter_002:rsp_src_valid -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_002_rsp_src_startofpacket                                                                   : std_logic;                      -- limiter_002:rsp_src_startofpacket -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_002_rsp_src_data                                                                            : std_logic_vector(126 downto 0); -- limiter_002:rsp_src_data -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_002_rsp_src_channel                                                                         : std_logic_vector(11 downto 0);  -- limiter_002:rsp_src_channel -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_002_rsp_src_ready                                                                           : std_logic;                      -- mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                                   : std_logic;                      -- burst_adapter:source0_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                         : std_logic;                      -- burst_adapter:source0_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                 : std_logic;                      -- burst_adapter:source0_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                          : std_logic_vector(126 downto 0); -- burst_adapter:source0_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                         : std_logic;                      -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                       : std_logic_vector(11 downto 0);  -- burst_adapter:source0_channel -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_001:source0_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                     : std_logic;                      -- burst_adapter_001:source0_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_001:source0_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_001:source0_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                     : std_logic;                      -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_001:source0_channel -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_002_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_002:source0_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_002_source0_valid                                                                     : std_logic;                      -- burst_adapter_002:source0_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_002_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_002:source0_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_002_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_002:source0_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_002_source0_ready                                                                     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	signal burst_adapter_002_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_002:source0_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_003_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_003:source0_endofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_003_source0_valid                                                                     : std_logic;                      -- burst_adapter_003:source0_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_003_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_003:source0_startofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_003_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_003:source0_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_003_source0_ready                                                                     : std_logic;                      -- mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	signal burst_adapter_003_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_003:source0_channel -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_004_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_004:source0_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_004_source0_valid                                                                     : std_logic;                      -- burst_adapter_004:source0_valid -> button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_004_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_004:source0_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_004_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_004:source0_data -> button_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_004_source0_ready                                                                     : std_logic;                      -- button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	signal burst_adapter_004_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_004:source0_channel -> button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_005_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_005:source0_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_005_source0_valid                                                                     : std_logic;                      -- burst_adapter_005:source0_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_005_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_005:source0_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_005_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_005:source0_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_005_source0_ready                                                                     : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_005:source0_ready
	signal burst_adapter_005_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_005:source0_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_006_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_006:source0_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_006_source0_valid                                                                     : std_logic;                      -- burst_adapter_006:source0_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_006_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_006:source0_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_006_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_006:source0_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_006_source0_ready                                                                     : std_logic;                      -- timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_006:source0_ready
	signal burst_adapter_006_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_006:source0_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_007_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_007:source0_endofpacket -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_007_source0_valid                                                                     : std_logic;                      -- burst_adapter_007:source0_valid -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_007_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_007:source0_startofpacket -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_007_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_007:source0_data -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_007_source0_ready                                                                     : std_logic;                      -- spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_007:source0_ready
	signal burst_adapter_007_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_007:source0_channel -> spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_008_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_008:source0_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_008_source0_valid                                                                     : std_logic;                      -- burst_adapter_008:source0_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_008_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_008:source0_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_008_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_008:source0_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_008_source0_ready                                                                     : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_008:source0_ready
	signal burst_adapter_008_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_008:source0_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_009_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_009:source0_endofpacket -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_009_source0_valid                                                                     : std_logic;                      -- burst_adapter_009:source0_valid -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_009_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_009:source0_startofpacket -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_009_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_009:source0_data -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_009_source0_ready                                                                     : std_logic;                      -- spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_009:source0_ready
	signal burst_adapter_009_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_009:source0_channel -> spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_010_source0_endofpacket                                                               : std_logic;                      -- burst_adapter_010:source0_endofpacket -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_010_source0_valid                                                                     : std_logic;                      -- burst_adapter_010:source0_valid -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_010_source0_startofpacket                                                             : std_logic;                      -- burst_adapter_010:source0_startofpacket -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_010_source0_data                                                                      : std_logic_vector(126 downto 0); -- burst_adapter_010:source0_data -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_010_source0_ready                                                                     : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_010:source0_ready
	signal burst_adapter_010_source0_channel                                                                   : std_logic_vector(11 downto 0);  -- burst_adapter_010:source0_channel -> no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                      : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmv_master_interface_0_avalon_master_translator:reset, cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:in_reset, crosser_007:in_reset, crosser_008:in_reset, crosser_009:in_reset, crosser_010:in_reset, crosser_011:in_reset, crosser_012:in_reset, crosser_013:in_reset, crosser_014:in_reset, crosser_015:out_reset, crosser_016:out_reset, crosser_017:out_reset, crosser_018:out_reset, crosser_019:out_reset, crosser_020:out_reset, crosser_021:out_reset, crosser_022:out_reset, crosser_023:out_reset, crosser_024:out_reset, crosser_025:out_reset, crosser_026:out_reset, crosser_027:out_reset, crosser_028:out_reset, crosser_029:out_reset, dvi_master_interface_0_avalon_master_translator:reset, dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:reset, id_router:reset, id_router_001:reset, id_router_002:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, limiter_002:reset, mm_clock_crossing_bridge_io:m0_reset, mm_clock_crossing_bridge_io_m0_translator:reset, mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:reset, nios2_qsys_data_master_translator:reset, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_instruction_master_translator:reset, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_jtag_debug_module_translator:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory:reset, onchip_memory_s1_translator:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, rst_controller_reset_out_reset:in, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset]
	signal rst_controller_001_reset_out_reset                                                                  : std_logic;                      -- rst_controller_001:reset_out -> [burst_adapter_003:reset, burst_adapter_004:reset, burst_adapter_005:reset, burst_adapter_006:reset, burst_adapter_007:reset, burst_adapter_008:reset, burst_adapter_009:reset, burst_adapter_010:reset, button_s1_translator:reset, button_s1_translator_avalon_universal_slave_0_agent:reset, button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_011:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:out_reset, crosser_008:out_reset, crosser_009:out_reset, crosser_010:out_reset, crosser_011:out_reset, crosser_012:out_reset, crosser_013:out_reset, crosser_014:out_reset, crosser_015:in_reset, crosser_016:in_reset, crosser_017:in_reset, crosser_018:in_reset, crosser_019:in_reset, crosser_020:in_reset, crosser_021:in_reset, crosser_022:in_reset, crosser_023:in_reset, crosser_024:in_reset, crosser_025:in_reset, crosser_026:in_reset, crosser_027:in_reset, crosser_028:in_reset, crosser_029:in_reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_010:reset, id_router_011:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mm_clock_crossing_bridge_io:s0_reset, mm_clock_crossing_bridge_io_s0_translator:reset, mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:reset, mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, no_of_cam_channels_s1_translator:reset, no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent:reset, no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rst_controller_001_reset_out_reset:in, spi_1_spi_control_port_translator:reset, spi_1_spi_control_port_translator_avalon_universal_slave_0_agent:reset, spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, spi_2_spi_control_port_translator:reset, spi_2_spi_control_port_translator_avalon_universal_slave_0_agent:reset, spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal rst_controller_002_reset_out_reset                                                                  : std_logic;                      -- rst_controller_002:reset_out -> [cmd_xbar_mux_009:reset, id_router_009:reset, mem_if_ddr2_emif_avl_translator:reset, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:reset, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_009:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset]
	signal mem_if_ddr2_emif_afi_reset_reset                                                                    : std_logic;                      -- mem_if_ddr2_emif:afi_reset_n -> mem_if_ddr2_emif_afi_reset_reset:in
	signal cmd_xbar_demux_src0_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                            : std_logic_vector(126 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                         : std_logic_vector(11 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                           : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                            : std_logic_vector(126 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                         : std_logic_vector(11 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                           : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                       : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                       : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> burst_adapter_002:sink0_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> burst_adapter_002:sink0_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> burst_adapter_002:sink0_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src2_data -> burst_adapter_002:sink0_data
	signal cmd_xbar_demux_001_src2_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src2_channel -> burst_adapter_002:sink0_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                     : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                           : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                   : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                            : std_logic_vector(126 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                         : std_logic_vector(11 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                           : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                     : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                           : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                   : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                            : std_logic_vector(126 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                         : std_logic_vector(11 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                           : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                       : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal limiter_cmd_src_endofpacket                                                                         : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                       : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                                : std_logic_vector(126 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                             : std_logic_vector(11 downto 0);  -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                               : std_logic;                      -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                        : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                              : std_logic;                      -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                                      : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                               : std_logic_vector(126 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                            : std_logic_vector(11 downto 0);  -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                              : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal limiter_001_cmd_src_endofpacket                                                                     : std_logic;                      -- limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal limiter_001_cmd_src_startofpacket                                                                   : std_logic;                      -- limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal limiter_001_cmd_src_data                                                                            : std_logic_vector(126 downto 0); -- limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	signal limiter_001_cmd_src_channel                                                                         : std_logic_vector(11 downto 0);  -- limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	signal limiter_001_cmd_src_ready                                                                           : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                    : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                          : std_logic;                      -- rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                  : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                           : std_logic_vector(126 downto 0); -- rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	signal rsp_xbar_mux_001_src_channel                                                                        : std_logic_vector(11 downto 0);  -- rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	signal rsp_xbar_mux_001_src_ready                                                                          : std_logic;                      -- limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	signal limiter_002_cmd_src_endofpacket                                                                     : std_logic;                      -- limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	signal limiter_002_cmd_src_startofpacket                                                                   : std_logic;                      -- limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	signal limiter_002_cmd_src_data                                                                            : std_logic_vector(126 downto 0); -- limiter_002:cmd_src_data -> cmd_xbar_demux_002:sink_data
	signal limiter_002_cmd_src_channel                                                                         : std_logic_vector(11 downto 0);  -- limiter_002:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	signal limiter_002_cmd_src_ready                                                                           : std_logic;                      -- cmd_xbar_demux_002:sink_ready -> limiter_002:cmd_src_ready
	signal rsp_xbar_mux_002_src_endofpacket                                                                    : std_logic;                      -- rsp_xbar_mux_002:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	signal rsp_xbar_mux_002_src_valid                                                                          : std_logic;                      -- rsp_xbar_mux_002:src_valid -> limiter_002:rsp_sink_valid
	signal rsp_xbar_mux_002_src_startofpacket                                                                  : std_logic;                      -- rsp_xbar_mux_002:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	signal rsp_xbar_mux_002_src_data                                                                           : std_logic_vector(126 downto 0); -- rsp_xbar_mux_002:src_data -> limiter_002:rsp_sink_data
	signal rsp_xbar_mux_002_src_channel                                                                        : std_logic_vector(11 downto 0);  -- rsp_xbar_mux_002:src_channel -> limiter_002:rsp_sink_channel
	signal rsp_xbar_mux_002_src_ready                                                                          : std_logic;                      -- limiter_002:rsp_sink_ready -> rsp_xbar_mux_002:src_ready
	signal addr_router_003_src_endofpacket                                                                     : std_logic;                      -- addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	signal addr_router_003_src_valid                                                                           : std_logic;                      -- addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	signal addr_router_003_src_startofpacket                                                                   : std_logic;                      -- addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	signal addr_router_003_src_data                                                                            : std_logic_vector(126 downto 0); -- addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	signal addr_router_003_src_channel                                                                         : std_logic_vector(11 downto 0);  -- addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	signal addr_router_003_src_ready                                                                           : std_logic;                      -- cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	signal width_adapter_004_src_ready                                                                         : std_logic;                      -- dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_004:out_ready
	signal addr_router_004_src_endofpacket                                                                     : std_logic;                      -- addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	signal addr_router_004_src_valid                                                                           : std_logic;                      -- addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	signal addr_router_004_src_startofpacket                                                                   : std_logic;                      -- addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	signal addr_router_004_src_data                                                                            : std_logic_vector(234 downto 0); -- addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	signal addr_router_004_src_channel                                                                         : std_logic_vector(11 downto 0);  -- addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	signal addr_router_004_src_ready                                                                           : std_logic;                      -- cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	signal width_adapter_005_src_ready                                                                         : std_logic;                      -- cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_005:out_ready
	signal cmd_xbar_mux_src_endofpacket                                                                        : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> burst_adapter:sink0_endofpacket
	signal cmd_xbar_mux_src_valid                                                                              : std_logic;                      -- cmd_xbar_mux:src_valid -> burst_adapter:sink0_valid
	signal cmd_xbar_mux_src_startofpacket                                                                      : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> burst_adapter:sink0_startofpacket
	signal cmd_xbar_mux_src_data                                                                               : std_logic_vector(126 downto 0); -- cmd_xbar_mux:src_data -> burst_adapter:sink0_data
	signal cmd_xbar_mux_src_channel                                                                            : std_logic_vector(11 downto 0);  -- cmd_xbar_mux:src_channel -> burst_adapter:sink0_channel
	signal cmd_xbar_mux_src_ready                                                                              : std_logic;                      -- burst_adapter:sink0_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                           : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                 : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                         : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                  : std_logic_vector(126 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                               : std_logic_vector(11 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                 : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_001:src_valid -> burst_adapter_001:sink0_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_001:src_data -> burst_adapter_001:sink0_data
	signal cmd_xbar_mux_001_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_001:src_channel -> burst_adapter_001:sink0_channel
	signal cmd_xbar_mux_001_src_ready                                                                          : std_logic;                      -- burst_adapter_001:sink0_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                       : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                             : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                     : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_demux_001_src2_ready                                                                       : std_logic;                      -- burst_adapter_002:sink0_ready -> cmd_xbar_demux_001:src2_ready
	signal id_router_002_src_endofpacket                                                                       : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                             : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                     : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal crosser_out_ready                                                                                   : std_logic;                      -- burst_adapter_003:sink0_ready -> crosser:out_ready
	signal id_router_003_src_endofpacket                                                                       : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                             : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                     : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_004:src_endofpacket -> burst_adapter_004:sink0_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_004:src_valid -> burst_adapter_004:sink0_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_004:src_startofpacket -> burst_adapter_004:sink0_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_004:src_data -> burst_adapter_004:sink0_data
	signal cmd_xbar_mux_004_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_004:src_channel -> burst_adapter_004:sink0_channel
	signal cmd_xbar_mux_004_src_ready                                                                          : std_logic;                      -- burst_adapter_004:sink0_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                       : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                             : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                     : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_mux_005_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_005:src_endofpacket -> burst_adapter_005:sink0_endofpacket
	signal cmd_xbar_mux_005_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_005:src_valid -> burst_adapter_005:sink0_valid
	signal cmd_xbar_mux_005_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_005:src_startofpacket -> burst_adapter_005:sink0_startofpacket
	signal cmd_xbar_mux_005_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_005:src_data -> burst_adapter_005:sink0_data
	signal cmd_xbar_mux_005_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_005:src_channel -> burst_adapter_005:sink0_channel
	signal cmd_xbar_mux_005_src_ready                                                                          : std_logic;                      -- burst_adapter_005:sink0_ready -> cmd_xbar_mux_005:src_ready
	signal id_router_005_src_endofpacket                                                                       : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                             : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                     : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_mux_006_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_006:src_endofpacket -> burst_adapter_006:sink0_endofpacket
	signal cmd_xbar_mux_006_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_006:src_valid -> burst_adapter_006:sink0_valid
	signal cmd_xbar_mux_006_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_006:src_startofpacket -> burst_adapter_006:sink0_startofpacket
	signal cmd_xbar_mux_006_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_006:src_data -> burst_adapter_006:sink0_data
	signal cmd_xbar_mux_006_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_006:src_channel -> burst_adapter_006:sink0_channel
	signal cmd_xbar_mux_006_src_ready                                                                          : std_logic;                      -- burst_adapter_006:sink0_ready -> cmd_xbar_mux_006:src_ready
	signal id_router_006_src_endofpacket                                                                       : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                             : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                     : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_mux_007_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_007:src_endofpacket -> burst_adapter_007:sink0_endofpacket
	signal cmd_xbar_mux_007_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_007:src_valid -> burst_adapter_007:sink0_valid
	signal cmd_xbar_mux_007_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_007:src_startofpacket -> burst_adapter_007:sink0_startofpacket
	signal cmd_xbar_mux_007_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_007:src_data -> burst_adapter_007:sink0_data
	signal cmd_xbar_mux_007_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_007:src_channel -> burst_adapter_007:sink0_channel
	signal cmd_xbar_mux_007_src_ready                                                                          : std_logic;                      -- burst_adapter_007:sink0_ready -> cmd_xbar_mux_007:src_ready
	signal id_router_007_src_endofpacket                                                                       : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                             : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                     : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_mux_008_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_008:src_endofpacket -> burst_adapter_008:sink0_endofpacket
	signal cmd_xbar_mux_008_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_008:src_valid -> burst_adapter_008:sink0_valid
	signal cmd_xbar_mux_008_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_008:src_startofpacket -> burst_adapter_008:sink0_startofpacket
	signal cmd_xbar_mux_008_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_008:src_data -> burst_adapter_008:sink0_data
	signal cmd_xbar_mux_008_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_008:src_channel -> burst_adapter_008:sink0_channel
	signal cmd_xbar_mux_008_src_ready                                                                          : std_logic;                      -- burst_adapter_008:sink0_ready -> cmd_xbar_mux_008:src_ready
	signal id_router_008_src_endofpacket                                                                       : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                             : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                     : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_mux_009_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_009:src_endofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_009_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_009:src_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_009_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_009:src_startofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_009_src_data                                                                           : std_logic_vector(378 downto 0); -- cmd_xbar_mux_009:src_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_009_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_009:src_channel -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_009_src_ready                                                                          : std_logic;                      -- mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	signal id_router_009_src_endofpacket                                                                       : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                             : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                     : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                              : std_logic_vector(378 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_mux_010_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_010:src_endofpacket -> burst_adapter_009:sink0_endofpacket
	signal cmd_xbar_mux_010_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_010:src_valid -> burst_adapter_009:sink0_valid
	signal cmd_xbar_mux_010_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_010:src_startofpacket -> burst_adapter_009:sink0_startofpacket
	signal cmd_xbar_mux_010_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_010:src_data -> burst_adapter_009:sink0_data
	signal cmd_xbar_mux_010_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_010:src_channel -> burst_adapter_009:sink0_channel
	signal cmd_xbar_mux_010_src_ready                                                                          : std_logic;                      -- burst_adapter_009:sink0_ready -> cmd_xbar_mux_010:src_ready
	signal id_router_010_src_endofpacket                                                                       : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                             : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                     : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_mux_011_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_011:src_endofpacket -> burst_adapter_010:sink0_endofpacket
	signal cmd_xbar_mux_011_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_011:src_valid -> burst_adapter_010:sink0_valid
	signal cmd_xbar_mux_011_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_011:src_startofpacket -> burst_adapter_010:sink0_startofpacket
	signal cmd_xbar_mux_011_src_data                                                                           : std_logic_vector(126 downto 0); -- cmd_xbar_mux_011:src_data -> burst_adapter_010:sink0_data
	signal cmd_xbar_mux_011_src_channel                                                                        : std_logic_vector(11 downto 0);  -- cmd_xbar_mux_011:src_channel -> burst_adapter_010:sink0_channel
	signal cmd_xbar_mux_011_src_ready                                                                          : std_logic;                      -- burst_adapter_010:sink0_ready -> cmd_xbar_mux_011:src_ready
	signal id_router_011_src_endofpacket                                                                       : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                             : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                     : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                              : std_logic_vector(126 downto 0); -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                           : std_logic_vector(11 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_001_src9_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src9_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src9_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src9_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src9_data -> width_adapter:in_data
	signal cmd_xbar_demux_001_src9_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src9_channel -> width_adapter:in_channel
	signal cmd_xbar_demux_001_src9_ready                                                                       : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_demux_001:src9_ready
	signal width_adapter_src_endofpacket                                                                       : std_logic;                      -- width_adapter:out_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	signal width_adapter_src_valid                                                                             : std_logic;                      -- width_adapter:out_valid -> cmd_xbar_mux_009:sink0_valid
	signal width_adapter_src_startofpacket                                                                     : std_logic;                      -- width_adapter:out_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	signal width_adapter_src_data                                                                              : std_logic_vector(378 downto 0); -- width_adapter:out_data -> cmd_xbar_mux_009:sink0_data
	signal width_adapter_src_ready                                                                             : std_logic;                      -- cmd_xbar_mux_009:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                           : std_logic_vector(11 downto 0);  -- width_adapter:out_channel -> cmd_xbar_mux_009:sink0_channel
	signal cmd_xbar_demux_003_src0_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_003:src0_endofpacket -> width_adapter_001:in_endofpacket
	signal cmd_xbar_demux_003_src0_valid                                                                       : std_logic;                      -- cmd_xbar_demux_003:src0_valid -> width_adapter_001:in_valid
	signal cmd_xbar_demux_003_src0_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_003:src0_startofpacket -> width_adapter_001:in_startofpacket
	signal cmd_xbar_demux_003_src0_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_003:src0_data -> width_adapter_001:in_data
	signal cmd_xbar_demux_003_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_003:src0_channel -> width_adapter_001:in_channel
	signal cmd_xbar_demux_003_src0_ready                                                                       : std_logic;                      -- width_adapter_001:in_ready -> cmd_xbar_demux_003:src0_ready
	signal width_adapter_001_src_endofpacket                                                                   : std_logic;                      -- width_adapter_001:out_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	signal width_adapter_001_src_valid                                                                         : std_logic;                      -- width_adapter_001:out_valid -> cmd_xbar_mux_009:sink1_valid
	signal width_adapter_001_src_startofpacket                                                                 : std_logic;                      -- width_adapter_001:out_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	signal width_adapter_001_src_data                                                                          : std_logic_vector(378 downto 0); -- width_adapter_001:out_data -> cmd_xbar_mux_009:sink1_data
	signal width_adapter_001_src_ready                                                                         : std_logic;                      -- cmd_xbar_mux_009:sink1_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                       : std_logic_vector(11 downto 0);  -- width_adapter_001:out_channel -> cmd_xbar_mux_009:sink1_channel
	signal cmd_xbar_demux_004_src0_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_004:src0_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_demux_004_src0_valid                                                                       : std_logic;                      -- cmd_xbar_demux_004:src0_valid -> width_adapter_002:in_valid
	signal cmd_xbar_demux_004_src0_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src0_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_demux_004_src0_data                                                                        : std_logic_vector(234 downto 0); -- cmd_xbar_demux_004:src0_data -> width_adapter_002:in_data
	signal cmd_xbar_demux_004_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_004:src0_channel -> width_adapter_002:in_channel
	signal cmd_xbar_demux_004_src0_ready                                                                       : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_demux_004:src0_ready
	signal width_adapter_002_src_endofpacket                                                                   : std_logic;                      -- width_adapter_002:out_endofpacket -> cmd_xbar_mux_009:sink2_endofpacket
	signal width_adapter_002_src_valid                                                                         : std_logic;                      -- width_adapter_002:out_valid -> cmd_xbar_mux_009:sink2_valid
	signal width_adapter_002_src_startofpacket                                                                 : std_logic;                      -- width_adapter_002:out_startofpacket -> cmd_xbar_mux_009:sink2_startofpacket
	signal width_adapter_002_src_data                                                                          : std_logic_vector(378 downto 0); -- width_adapter_002:out_data -> cmd_xbar_mux_009:sink2_data
	signal width_adapter_002_src_ready                                                                         : std_logic;                      -- cmd_xbar_mux_009:sink2_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                       : std_logic_vector(11 downto 0);  -- width_adapter_002:out_channel -> cmd_xbar_mux_009:sink2_channel
	signal rsp_xbar_demux_009_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> width_adapter_003:in_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> width_adapter_003:in_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> width_adapter_003:in_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                        : std_logic_vector(378 downto 0); -- rsp_xbar_demux_009:src0_data -> width_adapter_003:in_data
	signal rsp_xbar_demux_009_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_009:src0_channel -> width_adapter_003:in_channel
	signal rsp_xbar_demux_009_src0_ready                                                                       : std_logic;                      -- width_adapter_003:in_ready -> rsp_xbar_demux_009:src0_ready
	signal width_adapter_003_src_endofpacket                                                                   : std_logic;                      -- width_adapter_003:out_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal width_adapter_003_src_valid                                                                         : std_logic;                      -- width_adapter_003:out_valid -> rsp_xbar_mux_001:sink9_valid
	signal width_adapter_003_src_startofpacket                                                                 : std_logic;                      -- width_adapter_003:out_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal width_adapter_003_src_data                                                                          : std_logic_vector(126 downto 0); -- width_adapter_003:out_data -> rsp_xbar_mux_001:sink9_data
	signal width_adapter_003_src_ready                                                                         : std_logic;                      -- rsp_xbar_mux_001:sink9_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                       : std_logic_vector(11 downto 0);  -- width_adapter_003:out_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_009:src1_endofpacket -> width_adapter_004:in_endofpacket
	signal rsp_xbar_demux_009_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_009:src1_valid -> width_adapter_004:in_valid
	signal rsp_xbar_demux_009_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_009:src1_startofpacket -> width_adapter_004:in_startofpacket
	signal rsp_xbar_demux_009_src1_data                                                                        : std_logic_vector(378 downto 0); -- rsp_xbar_demux_009:src1_data -> width_adapter_004:in_data
	signal rsp_xbar_demux_009_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_009:src1_channel -> width_adapter_004:in_channel
	signal rsp_xbar_demux_009_src1_ready                                                                       : std_logic;                      -- width_adapter_004:in_ready -> rsp_xbar_demux_009:src1_ready
	signal width_adapter_004_src_endofpacket                                                                   : std_logic;                      -- width_adapter_004:out_endofpacket -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal width_adapter_004_src_valid                                                                         : std_logic;                      -- width_adapter_004:out_valid -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	signal width_adapter_004_src_startofpacket                                                                 : std_logic;                      -- width_adapter_004:out_startofpacket -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal width_adapter_004_src_data                                                                          : std_logic_vector(126 downto 0); -- width_adapter_004:out_data -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	signal width_adapter_004_src_channel                                                                       : std_logic_vector(11 downto 0);  -- width_adapter_004:out_channel -> dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_009_src2_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_009:src2_endofpacket -> width_adapter_005:in_endofpacket
	signal rsp_xbar_demux_009_src2_valid                                                                       : std_logic;                      -- rsp_xbar_demux_009:src2_valid -> width_adapter_005:in_valid
	signal rsp_xbar_demux_009_src2_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_009:src2_startofpacket -> width_adapter_005:in_startofpacket
	signal rsp_xbar_demux_009_src2_data                                                                        : std_logic_vector(378 downto 0); -- rsp_xbar_demux_009:src2_data -> width_adapter_005:in_data
	signal rsp_xbar_demux_009_src2_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_009:src2_channel -> width_adapter_005:in_channel
	signal rsp_xbar_demux_009_src2_ready                                                                       : std_logic;                      -- width_adapter_005:in_ready -> rsp_xbar_demux_009:src2_ready
	signal width_adapter_005_src_endofpacket                                                                   : std_logic;                      -- width_adapter_005:out_endofpacket -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal width_adapter_005_src_valid                                                                         : std_logic;                      -- width_adapter_005:out_valid -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	signal width_adapter_005_src_startofpacket                                                                 : std_logic;                      -- width_adapter_005:out_startofpacket -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal width_adapter_005_src_data                                                                          : std_logic_vector(234 downto 0); -- width_adapter_005:out_data -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	signal width_adapter_005_src_channel                                                                       : std_logic_vector(11 downto 0);  -- width_adapter_005:out_channel -> cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	signal crosser_out_endofpacket                                                                             : std_logic;                      -- crosser:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	signal crosser_out_valid                                                                                   : std_logic;                      -- crosser:out_valid -> burst_adapter_003:sink0_valid
	signal crosser_out_startofpacket                                                                           : std_logic;                      -- crosser:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	signal crosser_out_data                                                                                    : std_logic_vector(126 downto 0); -- crosser:out_data -> burst_adapter_003:sink0_data
	signal crosser_out_channel                                                                                 : std_logic_vector(11 downto 0);  -- crosser:out_channel -> burst_adapter_003:sink0_channel
	signal cmd_xbar_demux_001_src3_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> crosser:in_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> crosser:in_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> crosser:in_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src3_data -> crosser:in_data
	signal cmd_xbar_demux_001_src3_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src3_channel -> crosser:in_channel
	signal cmd_xbar_demux_001_src3_ready                                                                       : std_logic;                      -- crosser:in_ready -> cmd_xbar_demux_001:src3_ready
	signal crosser_001_out_endofpacket                                                                         : std_logic;                      -- crosser_001:out_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal crosser_001_out_valid                                                                               : std_logic;                      -- crosser_001:out_valid -> cmd_xbar_mux_004:sink0_valid
	signal crosser_001_out_startofpacket                                                                       : std_logic;                      -- crosser_001:out_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal crosser_001_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_001:out_data -> cmd_xbar_mux_004:sink0_data
	signal crosser_001_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_001:out_channel -> cmd_xbar_mux_004:sink0_channel
	signal crosser_001_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_004:sink0_ready -> crosser_001:out_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> crosser_001:in_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> crosser_001:in_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> crosser_001:in_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src4_data -> crosser_001:in_data
	signal cmd_xbar_demux_001_src4_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src4_channel -> crosser_001:in_channel
	signal cmd_xbar_demux_001_src4_ready                                                                       : std_logic;                      -- crosser_001:in_ready -> cmd_xbar_demux_001:src4_ready
	signal crosser_002_out_endofpacket                                                                         : std_logic;                      -- crosser_002:out_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	signal crosser_002_out_valid                                                                               : std_logic;                      -- crosser_002:out_valid -> cmd_xbar_mux_005:sink0_valid
	signal crosser_002_out_startofpacket                                                                       : std_logic;                      -- crosser_002:out_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	signal crosser_002_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_002:out_data -> cmd_xbar_mux_005:sink0_data
	signal crosser_002_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_002:out_channel -> cmd_xbar_mux_005:sink0_channel
	signal crosser_002_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_005:sink0_ready -> crosser_002:out_ready
	signal cmd_xbar_demux_001_src5_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> crosser_002:in_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> crosser_002:in_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> crosser_002:in_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src5_data -> crosser_002:in_data
	signal cmd_xbar_demux_001_src5_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src5_channel -> crosser_002:in_channel
	signal cmd_xbar_demux_001_src5_ready                                                                       : std_logic;                      -- crosser_002:in_ready -> cmd_xbar_demux_001:src5_ready
	signal crosser_003_out_endofpacket                                                                         : std_logic;                      -- crosser_003:out_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	signal crosser_003_out_valid                                                                               : std_logic;                      -- crosser_003:out_valid -> cmd_xbar_mux_006:sink0_valid
	signal crosser_003_out_startofpacket                                                                       : std_logic;                      -- crosser_003:out_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	signal crosser_003_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_003:out_data -> cmd_xbar_mux_006:sink0_data
	signal crosser_003_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_003:out_channel -> cmd_xbar_mux_006:sink0_channel
	signal crosser_003_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_006:sink0_ready -> crosser_003:out_ready
	signal cmd_xbar_demux_001_src6_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> crosser_003:in_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> crosser_003:in_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> crosser_003:in_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src6_data -> crosser_003:in_data
	signal cmd_xbar_demux_001_src6_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src6_channel -> crosser_003:in_channel
	signal cmd_xbar_demux_001_src6_ready                                                                       : std_logic;                      -- crosser_003:in_ready -> cmd_xbar_demux_001:src6_ready
	signal crosser_004_out_endofpacket                                                                         : std_logic;                      -- crosser_004:out_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	signal crosser_004_out_valid                                                                               : std_logic;                      -- crosser_004:out_valid -> cmd_xbar_mux_007:sink0_valid
	signal crosser_004_out_startofpacket                                                                       : std_logic;                      -- crosser_004:out_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	signal crosser_004_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_004:out_data -> cmd_xbar_mux_007:sink0_data
	signal crosser_004_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_004:out_channel -> cmd_xbar_mux_007:sink0_channel
	signal crosser_004_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_007:sink0_ready -> crosser_004:out_ready
	signal cmd_xbar_demux_001_src7_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src7_endofpacket -> crosser_004:in_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src7_valid -> crosser_004:in_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src7_startofpacket -> crosser_004:in_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src7_data -> crosser_004:in_data
	signal cmd_xbar_demux_001_src7_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src7_channel -> crosser_004:in_channel
	signal cmd_xbar_demux_001_src7_ready                                                                       : std_logic;                      -- crosser_004:in_ready -> cmd_xbar_demux_001:src7_ready
	signal crosser_005_out_endofpacket                                                                         : std_logic;                      -- crosser_005:out_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	signal crosser_005_out_valid                                                                               : std_logic;                      -- crosser_005:out_valid -> cmd_xbar_mux_008:sink0_valid
	signal crosser_005_out_startofpacket                                                                       : std_logic;                      -- crosser_005:out_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	signal crosser_005_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_005:out_data -> cmd_xbar_mux_008:sink0_data
	signal crosser_005_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_005:out_channel -> cmd_xbar_mux_008:sink0_channel
	signal crosser_005_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_008:sink0_ready -> crosser_005:out_ready
	signal cmd_xbar_demux_001_src8_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src8_endofpacket -> crosser_005:in_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src8_valid -> crosser_005:in_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src8_startofpacket -> crosser_005:in_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src8_data -> crosser_005:in_data
	signal cmd_xbar_demux_001_src8_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src8_channel -> crosser_005:in_channel
	signal cmd_xbar_demux_001_src8_ready                                                                       : std_logic;                      -- crosser_005:in_ready -> cmd_xbar_demux_001:src8_ready
	signal crosser_006_out_endofpacket                                                                         : std_logic;                      -- crosser_006:out_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	signal crosser_006_out_valid                                                                               : std_logic;                      -- crosser_006:out_valid -> cmd_xbar_mux_010:sink0_valid
	signal crosser_006_out_startofpacket                                                                       : std_logic;                      -- crosser_006:out_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	signal crosser_006_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_006:out_data -> cmd_xbar_mux_010:sink0_data
	signal crosser_006_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_006:out_channel -> cmd_xbar_mux_010:sink0_channel
	signal crosser_006_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_010:sink0_ready -> crosser_006:out_ready
	signal cmd_xbar_demux_001_src10_endofpacket                                                                : std_logic;                      -- cmd_xbar_demux_001:src10_endofpacket -> crosser_006:in_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                                      : std_logic;                      -- cmd_xbar_demux_001:src10_valid -> crosser_006:in_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                              : std_logic;                      -- cmd_xbar_demux_001:src10_startofpacket -> crosser_006:in_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                       : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src10_data -> crosser_006:in_data
	signal cmd_xbar_demux_001_src10_channel                                                                    : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src10_channel -> crosser_006:in_channel
	signal cmd_xbar_demux_001_src10_ready                                                                      : std_logic;                      -- crosser_006:in_ready -> cmd_xbar_demux_001:src10_ready
	signal crosser_007_out_endofpacket                                                                         : std_logic;                      -- crosser_007:out_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	signal crosser_007_out_valid                                                                               : std_logic;                      -- crosser_007:out_valid -> cmd_xbar_mux_011:sink0_valid
	signal crosser_007_out_startofpacket                                                                       : std_logic;                      -- crosser_007:out_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	signal crosser_007_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_007:out_data -> cmd_xbar_mux_011:sink0_data
	signal crosser_007_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_007:out_channel -> cmd_xbar_mux_011:sink0_channel
	signal crosser_007_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_011:sink0_ready -> crosser_007:out_ready
	signal cmd_xbar_demux_001_src11_endofpacket                                                                : std_logic;                      -- cmd_xbar_demux_001:src11_endofpacket -> crosser_007:in_endofpacket
	signal cmd_xbar_demux_001_src11_valid                                                                      : std_logic;                      -- cmd_xbar_demux_001:src11_valid -> crosser_007:in_valid
	signal cmd_xbar_demux_001_src11_startofpacket                                                              : std_logic;                      -- cmd_xbar_demux_001:src11_startofpacket -> crosser_007:in_startofpacket
	signal cmd_xbar_demux_001_src11_data                                                                       : std_logic_vector(126 downto 0); -- cmd_xbar_demux_001:src11_data -> crosser_007:in_data
	signal cmd_xbar_demux_001_src11_channel                                                                    : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_001:src11_channel -> crosser_007:in_channel
	signal cmd_xbar_demux_001_src11_ready                                                                      : std_logic;                      -- crosser_007:in_ready -> cmd_xbar_demux_001:src11_ready
	signal crosser_008_out_endofpacket                                                                         : std_logic;                      -- crosser_008:out_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal crosser_008_out_valid                                                                               : std_logic;                      -- crosser_008:out_valid -> cmd_xbar_mux_004:sink1_valid
	signal crosser_008_out_startofpacket                                                                       : std_logic;                      -- crosser_008:out_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal crosser_008_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_008:out_data -> cmd_xbar_mux_004:sink1_data
	signal crosser_008_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_008:out_channel -> cmd_xbar_mux_004:sink1_channel
	signal crosser_008_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_004:sink1_ready -> crosser_008:out_ready
	signal cmd_xbar_demux_002_src0_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src0_endofpacket -> crosser_008:in_endofpacket
	signal cmd_xbar_demux_002_src0_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src0_valid -> crosser_008:in_valid
	signal cmd_xbar_demux_002_src0_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src0_startofpacket -> crosser_008:in_startofpacket
	signal cmd_xbar_demux_002_src0_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_002:src0_data -> crosser_008:in_data
	signal cmd_xbar_demux_002_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_002:src0_channel -> crosser_008:in_channel
	signal cmd_xbar_demux_002_src0_ready                                                                       : std_logic;                      -- crosser_008:in_ready -> cmd_xbar_demux_002:src0_ready
	signal crosser_009_out_endofpacket                                                                         : std_logic;                      -- crosser_009:out_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	signal crosser_009_out_valid                                                                               : std_logic;                      -- crosser_009:out_valid -> cmd_xbar_mux_005:sink1_valid
	signal crosser_009_out_startofpacket                                                                       : std_logic;                      -- crosser_009:out_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	signal crosser_009_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_009:out_data -> cmd_xbar_mux_005:sink1_data
	signal crosser_009_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_009:out_channel -> cmd_xbar_mux_005:sink1_channel
	signal crosser_009_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_005:sink1_ready -> crosser_009:out_ready
	signal cmd_xbar_demux_002_src1_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src1_endofpacket -> crosser_009:in_endofpacket
	signal cmd_xbar_demux_002_src1_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src1_valid -> crosser_009:in_valid
	signal cmd_xbar_demux_002_src1_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src1_startofpacket -> crosser_009:in_startofpacket
	signal cmd_xbar_demux_002_src1_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_002:src1_data -> crosser_009:in_data
	signal cmd_xbar_demux_002_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_002:src1_channel -> crosser_009:in_channel
	signal cmd_xbar_demux_002_src1_ready                                                                       : std_logic;                      -- crosser_009:in_ready -> cmd_xbar_demux_002:src1_ready
	signal crosser_010_out_endofpacket                                                                         : std_logic;                      -- crosser_010:out_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	signal crosser_010_out_valid                                                                               : std_logic;                      -- crosser_010:out_valid -> cmd_xbar_mux_006:sink1_valid
	signal crosser_010_out_startofpacket                                                                       : std_logic;                      -- crosser_010:out_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	signal crosser_010_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_010:out_data -> cmd_xbar_mux_006:sink1_data
	signal crosser_010_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_010:out_channel -> cmd_xbar_mux_006:sink1_channel
	signal crosser_010_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_006:sink1_ready -> crosser_010:out_ready
	signal cmd_xbar_demux_002_src2_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src2_endofpacket -> crosser_010:in_endofpacket
	signal cmd_xbar_demux_002_src2_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src2_valid -> crosser_010:in_valid
	signal cmd_xbar_demux_002_src2_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src2_startofpacket -> crosser_010:in_startofpacket
	signal cmd_xbar_demux_002_src2_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_002:src2_data -> crosser_010:in_data
	signal cmd_xbar_demux_002_src2_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_002:src2_channel -> crosser_010:in_channel
	signal cmd_xbar_demux_002_src2_ready                                                                       : std_logic;                      -- crosser_010:in_ready -> cmd_xbar_demux_002:src2_ready
	signal crosser_011_out_endofpacket                                                                         : std_logic;                      -- crosser_011:out_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	signal crosser_011_out_valid                                                                               : std_logic;                      -- crosser_011:out_valid -> cmd_xbar_mux_007:sink1_valid
	signal crosser_011_out_startofpacket                                                                       : std_logic;                      -- crosser_011:out_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	signal crosser_011_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_011:out_data -> cmd_xbar_mux_007:sink1_data
	signal crosser_011_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_011:out_channel -> cmd_xbar_mux_007:sink1_channel
	signal crosser_011_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_007:sink1_ready -> crosser_011:out_ready
	signal cmd_xbar_demux_002_src3_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src3_endofpacket -> crosser_011:in_endofpacket
	signal cmd_xbar_demux_002_src3_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src3_valid -> crosser_011:in_valid
	signal cmd_xbar_demux_002_src3_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src3_startofpacket -> crosser_011:in_startofpacket
	signal cmd_xbar_demux_002_src3_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_002:src3_data -> crosser_011:in_data
	signal cmd_xbar_demux_002_src3_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_002:src3_channel -> crosser_011:in_channel
	signal cmd_xbar_demux_002_src3_ready                                                                       : std_logic;                      -- crosser_011:in_ready -> cmd_xbar_demux_002:src3_ready
	signal crosser_012_out_endofpacket                                                                         : std_logic;                      -- crosser_012:out_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	signal crosser_012_out_valid                                                                               : std_logic;                      -- crosser_012:out_valid -> cmd_xbar_mux_008:sink1_valid
	signal crosser_012_out_startofpacket                                                                       : std_logic;                      -- crosser_012:out_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	signal crosser_012_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_012:out_data -> cmd_xbar_mux_008:sink1_data
	signal crosser_012_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_012:out_channel -> cmd_xbar_mux_008:sink1_channel
	signal crosser_012_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_008:sink1_ready -> crosser_012:out_ready
	signal cmd_xbar_demux_002_src4_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src4_endofpacket -> crosser_012:in_endofpacket
	signal cmd_xbar_demux_002_src4_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src4_valid -> crosser_012:in_valid
	signal cmd_xbar_demux_002_src4_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src4_startofpacket -> crosser_012:in_startofpacket
	signal cmd_xbar_demux_002_src4_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_002:src4_data -> crosser_012:in_data
	signal cmd_xbar_demux_002_src4_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_002:src4_channel -> crosser_012:in_channel
	signal cmd_xbar_demux_002_src4_ready                                                                       : std_logic;                      -- crosser_012:in_ready -> cmd_xbar_demux_002:src4_ready
	signal crosser_013_out_endofpacket                                                                         : std_logic;                      -- crosser_013:out_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	signal crosser_013_out_valid                                                                               : std_logic;                      -- crosser_013:out_valid -> cmd_xbar_mux_010:sink1_valid
	signal crosser_013_out_startofpacket                                                                       : std_logic;                      -- crosser_013:out_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	signal crosser_013_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_013:out_data -> cmd_xbar_mux_010:sink1_data
	signal crosser_013_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_013:out_channel -> cmd_xbar_mux_010:sink1_channel
	signal crosser_013_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_010:sink1_ready -> crosser_013:out_ready
	signal cmd_xbar_demux_002_src5_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src5_endofpacket -> crosser_013:in_endofpacket
	signal cmd_xbar_demux_002_src5_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src5_valid -> crosser_013:in_valid
	signal cmd_xbar_demux_002_src5_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src5_startofpacket -> crosser_013:in_startofpacket
	signal cmd_xbar_demux_002_src5_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_002:src5_data -> crosser_013:in_data
	signal cmd_xbar_demux_002_src5_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_002:src5_channel -> crosser_013:in_channel
	signal cmd_xbar_demux_002_src5_ready                                                                       : std_logic;                      -- crosser_013:in_ready -> cmd_xbar_demux_002:src5_ready
	signal crosser_014_out_endofpacket                                                                         : std_logic;                      -- crosser_014:out_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	signal crosser_014_out_valid                                                                               : std_logic;                      -- crosser_014:out_valid -> cmd_xbar_mux_011:sink1_valid
	signal crosser_014_out_startofpacket                                                                       : std_logic;                      -- crosser_014:out_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	signal crosser_014_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_014:out_data -> cmd_xbar_mux_011:sink1_data
	signal crosser_014_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_014:out_channel -> cmd_xbar_mux_011:sink1_channel
	signal crosser_014_out_ready                                                                               : std_logic;                      -- cmd_xbar_mux_011:sink1_ready -> crosser_014:out_ready
	signal cmd_xbar_demux_002_src6_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src6_endofpacket -> crosser_014:in_endofpacket
	signal cmd_xbar_demux_002_src6_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src6_valid -> crosser_014:in_valid
	signal cmd_xbar_demux_002_src6_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src6_startofpacket -> crosser_014:in_startofpacket
	signal cmd_xbar_demux_002_src6_data                                                                        : std_logic_vector(126 downto 0); -- cmd_xbar_demux_002:src6_data -> crosser_014:in_data
	signal cmd_xbar_demux_002_src6_channel                                                                     : std_logic_vector(11 downto 0);  -- cmd_xbar_demux_002:src6_channel -> crosser_014:in_channel
	signal cmd_xbar_demux_002_src6_ready                                                                       : std_logic;                      -- crosser_014:in_ready -> cmd_xbar_demux_002:src6_ready
	signal crosser_015_out_endofpacket                                                                         : std_logic;                      -- crosser_015:out_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal crosser_015_out_valid                                                                               : std_logic;                      -- crosser_015:out_valid -> rsp_xbar_mux_001:sink3_valid
	signal crosser_015_out_startofpacket                                                                       : std_logic;                      -- crosser_015:out_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal crosser_015_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_015:out_data -> rsp_xbar_mux_001:sink3_data
	signal crosser_015_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_015:out_channel -> rsp_xbar_mux_001:sink3_channel
	signal crosser_015_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> crosser_015:out_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> crosser_015:in_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> crosser_015:in_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> crosser_015:in_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_003:src0_data -> crosser_015:in_data
	signal rsp_xbar_demux_003_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_003:src0_channel -> crosser_015:in_channel
	signal rsp_xbar_demux_003_src0_ready                                                                       : std_logic;                      -- crosser_015:in_ready -> rsp_xbar_demux_003:src0_ready
	signal crosser_016_out_endofpacket                                                                         : std_logic;                      -- crosser_016:out_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal crosser_016_out_valid                                                                               : std_logic;                      -- crosser_016:out_valid -> rsp_xbar_mux_001:sink4_valid
	signal crosser_016_out_startofpacket                                                                       : std_logic;                      -- crosser_016:out_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal crosser_016_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_016:out_data -> rsp_xbar_mux_001:sink4_data
	signal crosser_016_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_016:out_channel -> rsp_xbar_mux_001:sink4_channel
	signal crosser_016_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> crosser_016:out_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> crosser_016:in_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> crosser_016:in_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> crosser_016:in_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_004:src0_data -> crosser_016:in_data
	signal rsp_xbar_demux_004_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_004:src0_channel -> crosser_016:in_channel
	signal rsp_xbar_demux_004_src0_ready                                                                       : std_logic;                      -- crosser_016:in_ready -> rsp_xbar_demux_004:src0_ready
	signal crosser_017_out_endofpacket                                                                         : std_logic;                      -- crosser_017:out_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	signal crosser_017_out_valid                                                                               : std_logic;                      -- crosser_017:out_valid -> rsp_xbar_mux_002:sink0_valid
	signal crosser_017_out_startofpacket                                                                       : std_logic;                      -- crosser_017:out_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	signal crosser_017_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_017:out_data -> rsp_xbar_mux_002:sink0_data
	signal crosser_017_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_017:out_channel -> rsp_xbar_mux_002:sink0_channel
	signal crosser_017_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink0_ready -> crosser_017:out_ready
	signal rsp_xbar_demux_004_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src1_endofpacket -> crosser_017:in_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_004:src1_valid -> crosser_017:in_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_004:src1_startofpacket -> crosser_017:in_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_004:src1_data -> crosser_017:in_data
	signal rsp_xbar_demux_004_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_004:src1_channel -> crosser_017:in_channel
	signal rsp_xbar_demux_004_src1_ready                                                                       : std_logic;                      -- crosser_017:in_ready -> rsp_xbar_demux_004:src1_ready
	signal crosser_018_out_endofpacket                                                                         : std_logic;                      -- crosser_018:out_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal crosser_018_out_valid                                                                               : std_logic;                      -- crosser_018:out_valid -> rsp_xbar_mux_001:sink5_valid
	signal crosser_018_out_startofpacket                                                                       : std_logic;                      -- crosser_018:out_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal crosser_018_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_018:out_data -> rsp_xbar_mux_001:sink5_data
	signal crosser_018_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_018:out_channel -> rsp_xbar_mux_001:sink5_channel
	signal crosser_018_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> crosser_018:out_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> crosser_018:in_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> crosser_018:in_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> crosser_018:in_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_005:src0_data -> crosser_018:in_data
	signal rsp_xbar_demux_005_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_005:src0_channel -> crosser_018:in_channel
	signal rsp_xbar_demux_005_src0_ready                                                                       : std_logic;                      -- crosser_018:in_ready -> rsp_xbar_demux_005:src0_ready
	signal crosser_019_out_endofpacket                                                                         : std_logic;                      -- crosser_019:out_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	signal crosser_019_out_valid                                                                               : std_logic;                      -- crosser_019:out_valid -> rsp_xbar_mux_002:sink1_valid
	signal crosser_019_out_startofpacket                                                                       : std_logic;                      -- crosser_019:out_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	signal crosser_019_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_019:out_data -> rsp_xbar_mux_002:sink1_data
	signal crosser_019_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_019:out_channel -> rsp_xbar_mux_002:sink1_channel
	signal crosser_019_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink1_ready -> crosser_019:out_ready
	signal rsp_xbar_demux_005_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src1_endofpacket -> crosser_019:in_endofpacket
	signal rsp_xbar_demux_005_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_005:src1_valid -> crosser_019:in_valid
	signal rsp_xbar_demux_005_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_005:src1_startofpacket -> crosser_019:in_startofpacket
	signal rsp_xbar_demux_005_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_005:src1_data -> crosser_019:in_data
	signal rsp_xbar_demux_005_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_005:src1_channel -> crosser_019:in_channel
	signal rsp_xbar_demux_005_src1_ready                                                                       : std_logic;                      -- crosser_019:in_ready -> rsp_xbar_demux_005:src1_ready
	signal crosser_020_out_endofpacket                                                                         : std_logic;                      -- crosser_020:out_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal crosser_020_out_valid                                                                               : std_logic;                      -- crosser_020:out_valid -> rsp_xbar_mux_001:sink6_valid
	signal crosser_020_out_startofpacket                                                                       : std_logic;                      -- crosser_020:out_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal crosser_020_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_020:out_data -> rsp_xbar_mux_001:sink6_data
	signal crosser_020_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_020:out_channel -> rsp_xbar_mux_001:sink6_channel
	signal crosser_020_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> crosser_020:out_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> crosser_020:in_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> crosser_020:in_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> crosser_020:in_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_006:src0_data -> crosser_020:in_data
	signal rsp_xbar_demux_006_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_006:src0_channel -> crosser_020:in_channel
	signal rsp_xbar_demux_006_src0_ready                                                                       : std_logic;                      -- crosser_020:in_ready -> rsp_xbar_demux_006:src0_ready
	signal crosser_021_out_endofpacket                                                                         : std_logic;                      -- crosser_021:out_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	signal crosser_021_out_valid                                                                               : std_logic;                      -- crosser_021:out_valid -> rsp_xbar_mux_002:sink2_valid
	signal crosser_021_out_startofpacket                                                                       : std_logic;                      -- crosser_021:out_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	signal crosser_021_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_021:out_data -> rsp_xbar_mux_002:sink2_data
	signal crosser_021_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_021:out_channel -> rsp_xbar_mux_002:sink2_channel
	signal crosser_021_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink2_ready -> crosser_021:out_ready
	signal rsp_xbar_demux_006_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_006:src1_endofpacket -> crosser_021:in_endofpacket
	signal rsp_xbar_demux_006_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_006:src1_valid -> crosser_021:in_valid
	signal rsp_xbar_demux_006_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_006:src1_startofpacket -> crosser_021:in_startofpacket
	signal rsp_xbar_demux_006_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_006:src1_data -> crosser_021:in_data
	signal rsp_xbar_demux_006_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_006:src1_channel -> crosser_021:in_channel
	signal rsp_xbar_demux_006_src1_ready                                                                       : std_logic;                      -- crosser_021:in_ready -> rsp_xbar_demux_006:src1_ready
	signal crosser_022_out_endofpacket                                                                         : std_logic;                      -- crosser_022:out_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal crosser_022_out_valid                                                                               : std_logic;                      -- crosser_022:out_valid -> rsp_xbar_mux_001:sink7_valid
	signal crosser_022_out_startofpacket                                                                       : std_logic;                      -- crosser_022:out_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal crosser_022_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_022:out_data -> rsp_xbar_mux_001:sink7_data
	signal crosser_022_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_022:out_channel -> rsp_xbar_mux_001:sink7_channel
	signal crosser_022_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink7_ready -> crosser_022:out_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> crosser_022:in_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> crosser_022:in_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> crosser_022:in_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_007:src0_data -> crosser_022:in_data
	signal rsp_xbar_demux_007_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_007:src0_channel -> crosser_022:in_channel
	signal rsp_xbar_demux_007_src0_ready                                                                       : std_logic;                      -- crosser_022:in_ready -> rsp_xbar_demux_007:src0_ready
	signal crosser_023_out_endofpacket                                                                         : std_logic;                      -- crosser_023:out_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	signal crosser_023_out_valid                                                                               : std_logic;                      -- crosser_023:out_valid -> rsp_xbar_mux_002:sink3_valid
	signal crosser_023_out_startofpacket                                                                       : std_logic;                      -- crosser_023:out_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	signal crosser_023_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_023:out_data -> rsp_xbar_mux_002:sink3_data
	signal crosser_023_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_023:out_channel -> rsp_xbar_mux_002:sink3_channel
	signal crosser_023_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink3_ready -> crosser_023:out_ready
	signal rsp_xbar_demux_007_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_007:src1_endofpacket -> crosser_023:in_endofpacket
	signal rsp_xbar_demux_007_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_007:src1_valid -> crosser_023:in_valid
	signal rsp_xbar_demux_007_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_007:src1_startofpacket -> crosser_023:in_startofpacket
	signal rsp_xbar_demux_007_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_007:src1_data -> crosser_023:in_data
	signal rsp_xbar_demux_007_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_007:src1_channel -> crosser_023:in_channel
	signal rsp_xbar_demux_007_src1_ready                                                                       : std_logic;                      -- crosser_023:in_ready -> rsp_xbar_demux_007:src1_ready
	signal crosser_024_out_endofpacket                                                                         : std_logic;                      -- crosser_024:out_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal crosser_024_out_valid                                                                               : std_logic;                      -- crosser_024:out_valid -> rsp_xbar_mux_001:sink8_valid
	signal crosser_024_out_startofpacket                                                                       : std_logic;                      -- crosser_024:out_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal crosser_024_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_024:out_data -> rsp_xbar_mux_001:sink8_data
	signal crosser_024_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_024:out_channel -> rsp_xbar_mux_001:sink8_channel
	signal crosser_024_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink8_ready -> crosser_024:out_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> crosser_024:in_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> crosser_024:in_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> crosser_024:in_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_008:src0_data -> crosser_024:in_data
	signal rsp_xbar_demux_008_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_008:src0_channel -> crosser_024:in_channel
	signal rsp_xbar_demux_008_src0_ready                                                                       : std_logic;                      -- crosser_024:in_ready -> rsp_xbar_demux_008:src0_ready
	signal crosser_025_out_endofpacket                                                                         : std_logic;                      -- crosser_025:out_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	signal crosser_025_out_valid                                                                               : std_logic;                      -- crosser_025:out_valid -> rsp_xbar_mux_002:sink4_valid
	signal crosser_025_out_startofpacket                                                                       : std_logic;                      -- crosser_025:out_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	signal crosser_025_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_025:out_data -> rsp_xbar_mux_002:sink4_data
	signal crosser_025_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_025:out_channel -> rsp_xbar_mux_002:sink4_channel
	signal crosser_025_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink4_ready -> crosser_025:out_ready
	signal rsp_xbar_demux_008_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_008:src1_endofpacket -> crosser_025:in_endofpacket
	signal rsp_xbar_demux_008_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_008:src1_valid -> crosser_025:in_valid
	signal rsp_xbar_demux_008_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_008:src1_startofpacket -> crosser_025:in_startofpacket
	signal rsp_xbar_demux_008_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_008:src1_data -> crosser_025:in_data
	signal rsp_xbar_demux_008_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_008:src1_channel -> crosser_025:in_channel
	signal rsp_xbar_demux_008_src1_ready                                                                       : std_logic;                      -- crosser_025:in_ready -> rsp_xbar_demux_008:src1_ready
	signal crosser_026_out_endofpacket                                                                         : std_logic;                      -- crosser_026:out_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal crosser_026_out_valid                                                                               : std_logic;                      -- crosser_026:out_valid -> rsp_xbar_mux_001:sink10_valid
	signal crosser_026_out_startofpacket                                                                       : std_logic;                      -- crosser_026:out_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal crosser_026_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_026:out_data -> rsp_xbar_mux_001:sink10_data
	signal crosser_026_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_026:out_channel -> rsp_xbar_mux_001:sink10_channel
	signal crosser_026_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink10_ready -> crosser_026:out_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> crosser_026:in_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> crosser_026:in_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> crosser_026:in_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_010:src0_data -> crosser_026:in_data
	signal rsp_xbar_demux_010_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_010:src0_channel -> crosser_026:in_channel
	signal rsp_xbar_demux_010_src0_ready                                                                       : std_logic;                      -- crosser_026:in_ready -> rsp_xbar_demux_010:src0_ready
	signal crosser_027_out_endofpacket                                                                         : std_logic;                      -- crosser_027:out_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	signal crosser_027_out_valid                                                                               : std_logic;                      -- crosser_027:out_valid -> rsp_xbar_mux_002:sink5_valid
	signal crosser_027_out_startofpacket                                                                       : std_logic;                      -- crosser_027:out_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	signal crosser_027_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_027:out_data -> rsp_xbar_mux_002:sink5_data
	signal crosser_027_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_027:out_channel -> rsp_xbar_mux_002:sink5_channel
	signal crosser_027_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink5_ready -> crosser_027:out_ready
	signal rsp_xbar_demux_010_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_010:src1_endofpacket -> crosser_027:in_endofpacket
	signal rsp_xbar_demux_010_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_010:src1_valid -> crosser_027:in_valid
	signal rsp_xbar_demux_010_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_010:src1_startofpacket -> crosser_027:in_startofpacket
	signal rsp_xbar_demux_010_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_010:src1_data -> crosser_027:in_data
	signal rsp_xbar_demux_010_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_010:src1_channel -> crosser_027:in_channel
	signal rsp_xbar_demux_010_src1_ready                                                                       : std_logic;                      -- crosser_027:in_ready -> rsp_xbar_demux_010:src1_ready
	signal crosser_028_out_endofpacket                                                                         : std_logic;                      -- crosser_028:out_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	signal crosser_028_out_valid                                                                               : std_logic;                      -- crosser_028:out_valid -> rsp_xbar_mux_001:sink11_valid
	signal crosser_028_out_startofpacket                                                                       : std_logic;                      -- crosser_028:out_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	signal crosser_028_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_028:out_data -> rsp_xbar_mux_001:sink11_data
	signal crosser_028_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_028:out_channel -> rsp_xbar_mux_001:sink11_channel
	signal crosser_028_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_001:sink11_ready -> crosser_028:out_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> crosser_028:in_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> crosser_028:in_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> crosser_028:in_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_011:src0_data -> crosser_028:in_data
	signal rsp_xbar_demux_011_src0_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_011:src0_channel -> crosser_028:in_channel
	signal rsp_xbar_demux_011_src0_ready                                                                       : std_logic;                      -- crosser_028:in_ready -> rsp_xbar_demux_011:src0_ready
	signal crosser_029_out_endofpacket                                                                         : std_logic;                      -- crosser_029:out_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	signal crosser_029_out_valid                                                                               : std_logic;                      -- crosser_029:out_valid -> rsp_xbar_mux_002:sink6_valid
	signal crosser_029_out_startofpacket                                                                       : std_logic;                      -- crosser_029:out_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	signal crosser_029_out_data                                                                                : std_logic_vector(126 downto 0); -- crosser_029:out_data -> rsp_xbar_mux_002:sink6_data
	signal crosser_029_out_channel                                                                             : std_logic_vector(11 downto 0);  -- crosser_029:out_channel -> rsp_xbar_mux_002:sink6_channel
	signal crosser_029_out_ready                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink6_ready -> crosser_029:out_ready
	signal rsp_xbar_demux_011_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_011:src1_endofpacket -> crosser_029:in_endofpacket
	signal rsp_xbar_demux_011_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_011:src1_valid -> crosser_029:in_valid
	signal rsp_xbar_demux_011_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_011:src1_startofpacket -> crosser_029:in_startofpacket
	signal rsp_xbar_demux_011_src1_data                                                                        : std_logic_vector(126 downto 0); -- rsp_xbar_demux_011:src1_data -> crosser_029:in_data
	signal rsp_xbar_demux_011_src1_channel                                                                     : std_logic_vector(11 downto 0);  -- rsp_xbar_demux_011:src1_channel -> crosser_029:in_channel
	signal rsp_xbar_demux_011_src1_ready                                                                       : std_logic;                      -- crosser_029:in_ready -> rsp_xbar_demux_011:src1_ready
	signal limiter_cmd_valid_data                                                                              : std_logic_vector(11 downto 0);  -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal limiter_001_cmd_valid_data                                                                          : std_logic_vector(11 downto 0);  -- limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	signal limiter_002_cmd_valid_data                                                                          : std_logic_vector(11 downto 0);  -- limiter_002:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	signal irq_mapper_receiver0_irq                                                                            : std_logic;                      -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal nios2_qsys_d_irq_irq                                                                                : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_qsys:d_irq
	signal irq_mapper_receiver1_irq                                                                            : std_logic;                      -- irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_receiver_irq                                                                       : std_logic_vector(0 downto 0);   -- timer:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver2_irq                                                                            : std_logic;                      -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_001_receiver_irq                                                                   : std_logic_vector(0 downto 0);   -- spi_2:irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver3_irq                                                                            : std_logic;                      -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	signal irq_synchronizer_002_receiver_irq                                                                   : std_logic_vector(0 downto 0);   -- spi_1:irq -> irq_synchronizer_002:receiver_irq
	signal reset_reset_n_ports_inv                                                                             : std_logic;                      -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                           : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart:av_read_n
	signal led_s1_translator_avalon_anti_slave_0_write_ports_inv                                               : std_logic;                      -- led_s1_translator_avalon_anti_slave_0_write:inv -> led:write_n
	signal timer_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                      -- timer_s1_translator_avalon_anti_slave_0_write:inv -> timer:write_n
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv                               : std_logic;                      -- spi_2_spi_control_port_translator_avalon_anti_slave_0_write:inv -> spi_2:write_n
	signal spi_2_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv                                : std_logic;                      -- spi_2_spi_control_port_translator_avalon_anti_slave_0_read:inv -> spi_2:read_n
	signal mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_inv                                             : std_logic;                      -- mem_if_ddr2_emif_avl_waitrequest:inv -> mem_if_ddr2_emif_avl_translator:av_waitrequest
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv                               : std_logic;                      -- spi_1_spi_control_port_translator_avalon_anti_slave_0_write:inv -> spi_1:write_n
	signal spi_1_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv                                : std_logic;                      -- spi_1_spi_control_port_translator_avalon_anti_slave_0_read:inv -> spi_1:read_n
	signal no_of_cam_channels_s1_translator_avalon_anti_slave_0_write_ports_inv                                : std_logic;                      -- no_of_cam_channels_s1_translator_avalon_anti_slave_0_write:inv -> no_of_cam_channels:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                            : std_logic;                      -- rst_controller_reset_out_reset:inv -> [cmv_master_interface_0:RstxRBI, dvi_master_interface_0:RstxRBI, jtag_uart:rst_n, nios2_qsys:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                                        : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [button:reset_n, led:reset_n, no_of_cam_channels:reset_n, spi_1:reset_n, spi_2:reset_n, sysid:reset_n, timer:reset_n]
	signal mem_if_ddr2_emif_afi_reset_reset_ports_inv                                                          : std_logic;                      -- mem_if_ddr2_emif_afi_reset_reset:inv -> rst_controller_002:reset_in0

begin

	onchip_memory : component DE4_QSYS_onchip_memory
		port map (
			clk        => mem_if_ddr2_emif_afi_clk_clk,                               --   clk1.clk
			address    => onchip_memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			chipselect => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			clken      => onchip_memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			readdata   => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			write      => onchip_memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			writedata  => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset                              -- reset1.reset
		);

	mem_if_ddr2_emif : component DE4_QSYS_mem_if_ddr2_emif
		port map (
			pll_ref_clk       => clk_clk,                                                                --  pll_ref_clk.clk
			global_reset_n    => reset_reset_n,                                                          -- global_reset.reset_n
			soft_reset_n      => reset_reset_n,                                                          --   soft_reset.reset_n
			afi_clk           => mem_if_ddr2_emif_afi_clk_clk,                                           --      afi_clk.clk
			afi_half_clk      => open,                                                                   -- afi_half_clk.clk
			afi_reset_n       => mem_if_ddr2_emif_afi_reset_reset,                                       --    afi_reset.reset_n
			mem_a             => memory_mem_a,                                                           --       memory.mem_a
			mem_ba            => memory_mem_ba,                                                          --             .mem_ba
			mem_ck            => memory_mem_ck,                                                          --             .mem_ck
			mem_ck_n          => memory_mem_ck_n,                                                        --             .mem_ck_n
			mem_cke           => memory_mem_cke,                                                         --             .mem_cke
			mem_cs_n          => memory_mem_cs_n,                                                        --             .mem_cs_n
			mem_dm            => memory_mem_dm,                                                          --             .mem_dm
			mem_ras_n         => memory_mem_ras_n,                                                       --             .mem_ras_n
			mem_cas_n         => memory_mem_cas_n,                                                       --             .mem_cas_n
			mem_we_n          => memory_mem_we_n,                                                        --             .mem_we_n
			mem_dq            => memory_mem_dq,                                                          --             .mem_dq
			mem_dqs           => memory_mem_dqs,                                                         --             .mem_dqs
			mem_dqs_n         => memory_mem_dqs_n,                                                       --             .mem_dqs_n
			mem_odt           => memory_mem_odt,                                                         --             .mem_odt
			avl_ready         => mem_if_ddr2_emif_avl_waitrequest,                                       --          avl.waitrequest_n
			avl_burstbegin    => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_beginbursttransfer, --             .beginbursttransfer
			avl_addr          => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_address,            --             .address
			avl_rdata_valid   => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdatavalid,      --             .readdatavalid
			avl_rdata         => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdata,           --             .readdata
			avl_wdata         => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_writedata,          --             .writedata
			avl_be            => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_byteenable,         --             .byteenable
			avl_read_req      => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_read,               --             .read
			avl_write_req     => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_write,              --             .write
			avl_size          => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_burstcount,         --             .burstcount
			local_init_done   => open,                                                                   --       status.local_init_done
			local_cal_success => open,                                                                   --             .local_cal_success
			local_cal_fail    => open,                                                                   --             .local_cal_fail
			oct_rdn           => oct_rdn,                                                                --          oct.rdn
			oct_rup           => oct_rup                                                                 --             .rup
		);

	nios2_qsys : component DE4_QSYS_nios2_qsys
		port map (
			clk                                   => mem_if_ddr2_emif_afi_clk_clk,                                              --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                                  --                   reset_n.reset_n
			d_address                             => nios2_qsys_data_master_address,                                            --               data_master.address
			d_byteenable                          => nios2_qsys_data_master_byteenable,                                         --                          .byteenable
			d_read                                => nios2_qsys_data_master_read,                                               --                          .read
			d_readdata                            => nios2_qsys_data_master_readdata,                                           --                          .readdata
			d_waitrequest                         => nios2_qsys_data_master_waitrequest,                                        --                          .waitrequest
			d_write                               => nios2_qsys_data_master_write,                                              --                          .write
			d_writedata                           => nios2_qsys_data_master_writedata,                                          --                          .writedata
			d_burstcount                          => nios2_qsys_data_master_burstcount,                                         --                          .burstcount
			d_readdatavalid                       => nios2_qsys_data_master_readdatavalid,                                      --                          .readdatavalid
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_data_master_debugaccess,                                        --                          .debugaccess
			i_address                             => nios2_qsys_instruction_master_address,                                     --        instruction_master.address
			i_read                                => nios2_qsys_instruction_master_read,                                        --                          .read
			i_readdata                            => nios2_qsys_instruction_master_readdata,                                    --                          .readdata
			i_waitrequest                         => nios2_qsys_instruction_master_waitrequest,                                 --                          .waitrequest
			i_readdatavalid                       => nios2_qsys_instruction_master_readdatavalid,                               --                          .readdatavalid
			d_irq                                 => nios2_qsys_d_irq_irq,                                                      --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                                      --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address,       --         jtag_debug_module.address
			jtag_debug_module_begintransfer       => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer, --                          .begintransfer
			jtag_debug_module_byteenable          => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,    --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,   --                          .debugaccess
			jtag_debug_module_readdata            => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata,      --                          .readdata
			jtag_debug_module_select              => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect,    --                          .chipselect
			jtag_debug_module_write               => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write,         --                          .write
			jtag_debug_module_writedata           => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata,     --                          .writedata
			no_ci_readra                          => open                                                                       -- custom_instruction_master.readra
		);

	jtag_uart : component DE4_QSYS_jtag_uart
		port map (
			clk            => mem_if_ddr2_emif_afi_clk_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                   --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                    --               irq.irq
		);

	sysid : component DE4_QSYS_sysid
		port map (
			clock    => clk_clk,                                                       --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,                  --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	timer : component DE4_QSYS_timer
		port map (
			clk        => clk_clk,                                                 --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => timer_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_synchronizer_receiver_irq(0)                         --   irq.irq
		);

	led : component DE4_QSYS_led
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => led_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => led_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => led_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => led_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => led_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => led_export                                             -- external_connection.export
		);

	button : component DE4_QSYS_button
		port map (
			clk      => clk_clk,                                           --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => button_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => button_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => button_export                                      -- external_connection.export
		);

	mm_clock_crossing_bridge_io : component DE4_QSYS_mm_clock_crossing_bridge_io
		port map (
			m0_clk           => mem_if_ddr2_emif_afi_clk_clk,                                                --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,                                              -- m0_reset.reset
			s0_clk           => clk_clk,                                                                     --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset,                                          -- s0_reset.reset
			s0_waitrequest   => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdata,      --         .readdata
			s0_readdatavalid => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_burstcount,    --         .burstcount
			s0_writedata     => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_writedata,     --         .writedata
			s0_address       => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_address,       --         .address
			s0_write         => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_write,         --         .write
			s0_read          => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_read,          --         .read
			s0_byteenable    => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_debugaccess,   --         .debugaccess
			m0_waitrequest   => mm_clock_crossing_bridge_io_m0_waitrequest,                                  --       m0.waitrequest
			m0_readdata      => mm_clock_crossing_bridge_io_m0_readdata,                                     --         .readdata
			m0_readdatavalid => mm_clock_crossing_bridge_io_m0_readdatavalid,                                --         .readdatavalid
			m0_burstcount    => mm_clock_crossing_bridge_io_m0_burstcount,                                   --         .burstcount
			m0_writedata     => mm_clock_crossing_bridge_io_m0_writedata,                                    --         .writedata
			m0_address       => mm_clock_crossing_bridge_io_m0_address,                                      --         .address
			m0_write         => mm_clock_crossing_bridge_io_m0_write,                                        --         .write
			m0_read          => mm_clock_crossing_bridge_io_m0_read,                                         --         .read
			m0_byteenable    => mm_clock_crossing_bridge_io_m0_byteenable,                                   --         .byteenable
			m0_debugaccess   => mm_clock_crossing_bridge_io_m0_debugaccess                                   --         .debugaccess
		);

	spi_2 : component DE4_QSYS_spi_2
		port map (
			clk           => clk_clk,                                                               --              clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,                          --            reset.reset_n
			data_from_cpu => spi_2_spi_control_port_translator_avalon_anti_slave_0_writedata,       -- spi_control_port.writedata
			data_to_cpu   => spi_2_spi_control_port_translator_avalon_anti_slave_0_readdata,        --                 .readdata
			mem_addr      => spi_2_spi_control_port_translator_avalon_anti_slave_0_address,         --                 .address
			read_n        => spi_2_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv,  --                 .read_n
			spi_select    => spi_2_spi_control_port_translator_avalon_anti_slave_0_chipselect,      --                 .chipselect
			write_n       => spi_2_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv, --                 .write_n
			irq           => irq_synchronizer_001_receiver_irq(0),                                  --              irq.irq
			MISO          => spi_2_MISO,                                                            --         external.export
			MOSI          => spi_2_MOSI,                                                            --                 .export
			SCLK          => spi_2_SCLK,                                                            --                 .export
			SS_n          => spi_2_SS_n                                                             --                 .export
		);

	spi_1 : component DE4_QSYS_spi_2
		port map (
			clk           => clk_clk,                                                               --              clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,                          --            reset.reset_n
			data_from_cpu => spi_1_spi_control_port_translator_avalon_anti_slave_0_writedata,       -- spi_control_port.writedata
			data_to_cpu   => spi_1_spi_control_port_translator_avalon_anti_slave_0_readdata,        --                 .readdata
			mem_addr      => spi_1_spi_control_port_translator_avalon_anti_slave_0_address,         --                 .address
			read_n        => spi_1_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv,  --                 .read_n
			spi_select    => spi_1_spi_control_port_translator_avalon_anti_slave_0_chipselect,      --                 .chipselect
			write_n       => spi_1_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv, --                 .write_n
			irq           => irq_synchronizer_002_receiver_irq(0),                                  --              irq.irq
			MISO          => spi_1_MISO,                                                            --         external.export
			MOSI          => spi_1_MOSI,                                                            --                 .export
			SCLK          => spi_1_SCLK,                                                            --                 .export
			SS_n          => spi_1_SS_n                                                             --                 .export
		);

	no_of_cam_channels : component DE4_QSYS_no_of_cam_channels
		port map (
			clk        => clk_clk,                                                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                         --               reset.reset_n
			address    => no_of_cam_channels_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => no_of_cam_channels_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => no_of_cam_channels_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => no_of_cam_channels_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => no_of_cam_channels_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => no_of_cam_channels_export                                             -- external_connection.export
		);

	cmv_master_interface_0 : component DE4_QSYS_cmv_master_interface_0
		port map (
			ClkxCI          => mem_if_ddr2_emif_afi_clk_clk,                     --    clock_main.clk
			RstxRBI         => rst_controller_reset_out_reset_ports_inv,         --       reset_n.reset_n
			AMWritexSO      => cmv_master_interface_0_avalon_master_write,       -- avalon_master.write
			AMWriteDataxDO  => cmv_master_interface_0_avalon_master_writedata,   --              .writedata
			AMAddressxDO    => cmv_master_interface_0_avalon_master_address,     --              .address
			AMBurstCountxSO => cmv_master_interface_0_avalon_master_burstcount,  --              .burstcount
			AMWaitReqxSI    => cmv_master_interface_0_avalon_master_waitrequest, --              .waitrequest
			PixelValidxSI   => cmv_master_interface_PixelValidxSI,               --   conduit_end.export
			RowValidxSI     => cmv_master_interface_RowValidxSI,                 --              .export
			FrameValidxSI   => cmv_master_interface_FrameValidxSI,               --              .export
			DataInxDI       => cmv_master_interface_DataInxDI,                   --              .export
			ClkLvdsRxxCI    => cmv_master_interface_ClkLvdsRxxCI                 --              .export
		);

	dvi_master_interface_0 : component DE4_QSYS_dvi_master_interface_0
		port map (
			ClkxCI             => mem_if_ddr2_emif_afi_clk_clk,                       --    clock_main.clk
			RstxRBI            => rst_controller_reset_out_reset_ports_inv,           --       reset_n.reset_n
			AmWaitReqxSI       => dvi_master_interface_0_avalon_master_waitrequest,   -- avalon_master.waitrequest
			AmAddressxDO       => dvi_master_interface_0_avalon_master_address,       --              .address
			AmReadDataxDI      => dvi_master_interface_0_avalon_master_readdata,      --              .readdata
			AmReadxSO          => dvi_master_interface_0_avalon_master_read,          --              .read
			AmReadDataValidxSI => dvi_master_interface_0_avalon_master_readdatavalid, --              .readdatavalid
			AmBurstCountxDO    => dvi_master_interface_0_avalon_master_burstcount,    --              .burstcount
			ClkDvixCI          => dvi_master_interface_ClkDvixCI,                     --   conduit_end.export
			DviNewLinexDI      => dvi_master_interface_DviNewLinexDI,                 --              .export
			DviNewFramexDI     => dvi_master_interface_DviNewFramexDI,                --              .export
			DviPixelAvxSI      => dvi_master_interface_DviPixelAvxSI,                 --              .export
			DviDataOutxDO      => dvi_master_interface_DviDataOutxDO                  --              .export
		);

	nios2_qsys_instruction_master_translator : component DE4_QSYS_nios2_qsys_instruction_master_translator
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                     --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   --                     reset.reset
			uav_address       => nios2_qsys_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => nios2_qsys_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => nios2_qsys_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read           => nios2_qsys_instruction_master_read,                                               --                          .read
			av_readdata       => nios2_qsys_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid  => nios2_qsys_instruction_master_readdatavalid                                       --                          .readdatavalid
		);

	nios2_qsys_data_master_translator : component DE4_QSYS_nios2_qsys_data_master_translator
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                              --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address       => nios2_qsys_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => nios2_qsys_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => nios2_qsys_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => nios2_qsys_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => nios2_qsys_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => nios2_qsys_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => nios2_qsys_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => nios2_qsys_data_master_waitrequest,                                        --                          .waitrequest
			av_burstcount     => nios2_qsys_data_master_burstcount,                                         --                          .burstcount
			av_byteenable     => nios2_qsys_data_master_byteenable,                                         --                          .byteenable
			av_read           => nios2_qsys_data_master_read,                                               --                          .read
			av_readdata       => nios2_qsys_data_master_readdata,                                           --                          .readdata
			av_readdatavalid  => nios2_qsys_data_master_readdatavalid,                                      --                          .readdatavalid
			av_write          => nios2_qsys_data_master_write,                                              --                          .write
			av_writedata      => nios2_qsys_data_master_writedata,                                          --                          .writedata
			av_debugaccess    => nios2_qsys_data_master_debugaccess                                         --                          .debugaccess
		);

	mm_clock_crossing_bridge_io_m0_translator : component DE4_QSYS_mm_clock_crossing_bridge_io_m0_translator
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                      --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    --                     reset.reset
			uav_address       => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => mm_clock_crossing_bridge_io_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => mm_clock_crossing_bridge_io_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount     => mm_clock_crossing_bridge_io_m0_burstcount(0),                                      --                          .burstcount
			av_byteenable     => mm_clock_crossing_bridge_io_m0_byteenable,                                         --                          .byteenable
			av_read           => mm_clock_crossing_bridge_io_m0_read,                                               --                          .read
			av_readdata       => mm_clock_crossing_bridge_io_m0_readdata,                                           --                          .readdata
			av_readdatavalid  => mm_clock_crossing_bridge_io_m0_readdatavalid,                                      --                          .readdatavalid
			av_write          => mm_clock_crossing_bridge_io_m0_write,                                              --                          .write
			av_writedata      => mm_clock_crossing_bridge_io_m0_writedata,                                          --                          .writedata
			av_debugaccess    => mm_clock_crossing_bridge_io_m0_debugaccess                                         --                          .debugaccess
		);

	dvi_master_interface_0_avalon_master_translator : component DE4_QSYS_dvi_master_interface_0_avalon_master_translator
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                            --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                                          --                     reset.reset
			uav_address       => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => dvi_master_interface_0_avalon_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => dvi_master_interface_0_avalon_master_waitrequest,                                        --                          .waitrequest
			av_burstcount     => dvi_master_interface_0_avalon_master_burstcount,                                         --                          .burstcount
			av_read           => dvi_master_interface_0_avalon_master_read,                                               --                          .read
			av_readdata       => dvi_master_interface_0_avalon_master_readdata,                                           --                          .readdata
			av_readdatavalid  => dvi_master_interface_0_avalon_master_readdatavalid                                       --                          .readdatavalid
		);

	cmv_master_interface_0_avalon_master_translator : component DE4_QSYS_cmv_master_interface_0_avalon_master_translator
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                            --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                                          --                     reset.reset
			uav_address       => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => cmv_master_interface_0_avalon_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => cmv_master_interface_0_avalon_master_waitrequest,                                        --                          .waitrequest
			av_burstcount     => cmv_master_interface_0_avalon_master_burstcount,                                         --                          .burstcount
			av_write          => cmv_master_interface_0_avalon_master_write,                                              --                          .write
			av_writedata      => cmv_master_interface_0_avalon_master_writedata                                           --                          .writedata
		);

	nios2_qsys_jtag_debug_module_translator : component de4_qsys_nios2_qsys_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => mem_if_ddr2_emif_afi_clk_clk,                                                            --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                                          --                    reset.reset
			uav_address           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer      => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_byteenable         => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect         => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_debugaccess        => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_read               => open,                                                                                    --              (terminated)
			av_beginbursttransfer => open,                                                                                    --              (terminated)
			av_burstcount         => open,                                                                                    --              (terminated)
			av_readdatavalid      => '0',                                                                                     --              (terminated)
			av_waitrequest        => '0',                                                                                     --              (terminated)
			av_writebyteenable    => open,                                                                                    --              (terminated)
			av_lock               => open,                                                                                    --              (terminated)
			av_clken              => open,                                                                                    --              (terminated)
			uav_clken             => '0',                                                                                     --              (terminated)
			av_outputenable       => open                                                                                     --              (terminated)
		);

	onchip_memory_s1_translator : component de4_qsys_onchip_memory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 15,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => mem_if_ddr2_emif_afi_clk_clk,                                                --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => onchip_memory_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => onchip_memory_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable         => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect         => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken              => onchip_memory_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read               => open,                                                                        --              (terminated)
			av_begintransfer      => open,                                                                        --              (terminated)
			av_beginbursttransfer => open,                                                                        --              (terminated)
			av_burstcount         => open,                                                                        --              (terminated)
			av_readdatavalid      => '0',                                                                         --              (terminated)
			av_waitrequest        => '0',                                                                         --              (terminated)
			av_writebyteenable    => open,                                                                        --              (terminated)
			av_lock               => open,                                                                        --              (terminated)
			uav_clken             => '0',                                                                         --              (terminated)
			av_debugaccess        => open,                                                                        --              (terminated)
			av_outputenable       => open                                                                         --              (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator : component de4_qsys_jtag_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => mem_if_ddr2_emif_afi_clk_clk,                                                           --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest        => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect         => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer      => open,                                                                                   --              (terminated)
			av_beginbursttransfer => open,                                                                                   --              (terminated)
			av_burstcount         => open,                                                                                   --              (terminated)
			av_byteenable         => open,                                                                                   --              (terminated)
			av_readdatavalid      => '0',                                                                                    --              (terminated)
			av_writebyteenable    => open,                                                                                   --              (terminated)
			av_lock               => open,                                                                                   --              (terminated)
			av_clken              => open,                                                                                   --              (terminated)
			uav_clken             => '0',                                                                                    --              (terminated)
			av_debugaccess        => open,                                                                                   --              (terminated)
			av_outputenable       => open                                                                                    --              (terminated)
		);

	mm_clock_crossing_bridge_io_s0_translator : component de4_qsys_mm_clock_crossing_bridge_io_s0_translator
		generic map (
			AV_ADDRESS_W                   => 10,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                                                   --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                                        --                    reset.reset
			uav_address           => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount         => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable         => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid      => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest        => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess        => mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer      => open,                                                                                      --              (terminated)
			av_beginbursttransfer => open,                                                                                      --              (terminated)
			av_writebyteenable    => open,                                                                                      --              (terminated)
			av_lock               => open,                                                                                      --              (terminated)
			av_chipselect         => open,                                                                                      --              (terminated)
			av_clken              => open,                                                                                      --              (terminated)
			uav_clken             => '0',                                                                                       --              (terminated)
			av_outputenable       => open                                                                                       --              (terminated)
		);

	button_s1_translator : component de4_qsys_button_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                              --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                   --                    reset.reset
			uav_address           => button_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => button_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => button_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => button_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => button_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => button_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => button_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata           => button_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write              => open,                                                                 --              (terminated)
			av_read               => open,                                                                 --              (terminated)
			av_writedata          => open,                                                                 --              (terminated)
			av_begintransfer      => open,                                                                 --              (terminated)
			av_beginbursttransfer => open,                                                                 --              (terminated)
			av_burstcount         => open,                                                                 --              (terminated)
			av_byteenable         => open,                                                                 --              (terminated)
			av_readdatavalid      => '0',                                                                  --              (terminated)
			av_waitrequest        => '0',                                                                  --              (terminated)
			av_writebyteenable    => open,                                                                 --              (terminated)
			av_lock               => open,                                                                 --              (terminated)
			av_chipselect         => open,                                                                 --              (terminated)
			av_clken              => open,                                                                 --              (terminated)
			uav_clken             => '0',                                                                  --              (terminated)
			av_debugaccess        => open,                                                                 --              (terminated)
			av_outputenable       => open                                                                  --              (terminated)
		);

	led_s1_translator : component de4_qsys_button_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                           --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                --                    reset.reset
			uav_address           => led_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => led_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => led_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => led_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => led_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => led_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => led_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => led_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => led_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => led_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => led_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read               => open,                                                              --              (terminated)
			av_begintransfer      => open,                                                              --              (terminated)
			av_beginbursttransfer => open,                                                              --              (terminated)
			av_burstcount         => open,                                                              --              (terminated)
			av_byteenable         => open,                                                              --              (terminated)
			av_readdatavalid      => '0',                                                               --              (terminated)
			av_waitrequest        => '0',                                                               --              (terminated)
			av_writebyteenable    => open,                                                              --              (terminated)
			av_lock               => open,                                                              --              (terminated)
			av_clken              => open,                                                              --              (terminated)
			uav_clken             => '0',                                                               --              (terminated)
			av_debugaccess        => open,                                                              --              (terminated)
			av_outputenable       => open                                                               --              (terminated)
		);

	timer_s1_translator : component de4_qsys_timer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                             --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                  --                    reset.reset
			uav_address           => timer_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => timer_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => timer_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => timer_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => timer_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => timer_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => timer_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => timer_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read               => open,                                                                --              (terminated)
			av_begintransfer      => open,                                                                --              (terminated)
			av_beginbursttransfer => open,                                                                --              (terminated)
			av_burstcount         => open,                                                                --              (terminated)
			av_byteenable         => open,                                                                --              (terminated)
			av_readdatavalid      => '0',                                                                 --              (terminated)
			av_waitrequest        => '0',                                                                 --              (terminated)
			av_writebyteenable    => open,                                                                --              (terminated)
			av_lock               => open,                                                                --              (terminated)
			av_clken              => open,                                                                --              (terminated)
			uav_clken             => '0',                                                                 --              (terminated)
			av_debugaccess        => open,                                                                --              (terminated)
			av_outputenable       => open                                                                 --              (terminated)
		);

	spi_2_spi_control_port_translator : component de4_qsys_timer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                                           --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                                --                    reset.reset
			uav_address           => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => spi_2_spi_control_port_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => spi_2_spi_control_port_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => spi_2_spi_control_port_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => spi_2_spi_control_port_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => spi_2_spi_control_port_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => spi_2_spi_control_port_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer      => open,                                                                              --              (terminated)
			av_beginbursttransfer => open,                                                                              --              (terminated)
			av_burstcount         => open,                                                                              --              (terminated)
			av_byteenable         => open,                                                                              --              (terminated)
			av_readdatavalid      => '0',                                                                               --              (terminated)
			av_waitrequest        => '0',                                                                               --              (terminated)
			av_writebyteenable    => open,                                                                              --              (terminated)
			av_lock               => open,                                                                              --              (terminated)
			av_clken              => open,                                                                              --              (terminated)
			uav_clken             => '0',                                                                               --              (terminated)
			av_debugaccess        => open,                                                                              --              (terminated)
			av_outputenable       => open                                                                               --              (terminated)
		);

	sysid_control_slave_translator : component de4_qsys_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                                        --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                             --                    reset.reset
			uav_address           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata           => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write              => open,                                                                           --              (terminated)
			av_read               => open,                                                                           --              (terminated)
			av_writedata          => open,                                                                           --              (terminated)
			av_begintransfer      => open,                                                                           --              (terminated)
			av_beginbursttransfer => open,                                                                           --              (terminated)
			av_burstcount         => open,                                                                           --              (terminated)
			av_byteenable         => open,                                                                           --              (terminated)
			av_readdatavalid      => '0',                                                                            --              (terminated)
			av_waitrequest        => '0',                                                                            --              (terminated)
			av_writebyteenable    => open,                                                                           --              (terminated)
			av_lock               => open,                                                                           --              (terminated)
			av_chipselect         => open,                                                                           --              (terminated)
			av_clken              => open,                                                                           --              (terminated)
			uav_clken             => '0',                                                                            --              (terminated)
			av_debugaccess        => open,                                                                           --              (terminated)
			av_outputenable       => open                                                                            --              (terminated)
		);

	mem_if_ddr2_emif_avl_translator : component de4_qsys_mem_if_ddr2_emif_avl_translator
		generic map (
			AV_ADDRESS_W                   => 25,
			AV_DATA_W                      => 256,
			UAV_DATA_W                     => 256,
			AV_BURSTCOUNT_W                => 8,
			AV_BYTEENABLE_W                => 32,
			UAV_BYTEENABLE_W               => 32,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 13,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 32,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => mem_if_ddr2_emif_afi_clk_clk,                                                    --                      clk.clk
			reset                 => rst_controller_002_reset_out_reset,                                              --                    reset.reset
			uav_address           => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_beginbursttransfer => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_beginbursttransfer,          --                         .beginbursttransfer
			av_burstcount         => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable         => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid      => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest        => mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_inv,                         --                         .waitrequest
			av_begintransfer      => open,                                                                            --              (terminated)
			av_writebyteenable    => open,                                                                            --              (terminated)
			av_lock               => open,                                                                            --              (terminated)
			av_chipselect         => open,                                                                            --              (terminated)
			av_clken              => open,                                                                            --              (terminated)
			uav_clken             => '0',                                                                             --              (terminated)
			av_debugaccess        => open,                                                                            --              (terminated)
			av_outputenable       => open                                                                             --              (terminated)
		);

	spi_1_spi_control_port_translator : component de4_qsys_timer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                                           --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                                --                    reset.reset
			uav_address           => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => spi_1_spi_control_port_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => spi_1_spi_control_port_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => spi_1_spi_control_port_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => spi_1_spi_control_port_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => spi_1_spi_control_port_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => spi_1_spi_control_port_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer      => open,                                                                              --              (terminated)
			av_beginbursttransfer => open,                                                                              --              (terminated)
			av_burstcount         => open,                                                                              --              (terminated)
			av_byteenable         => open,                                                                              --              (terminated)
			av_readdatavalid      => '0',                                                                               --              (terminated)
			av_waitrequest        => '0',                                                                               --              (terminated)
			av_writebyteenable    => open,                                                                              --              (terminated)
			av_lock               => open,                                                                              --              (terminated)
			av_clken              => open,                                                                              --              (terminated)
			uav_clken             => '0',                                                                               --              (terminated)
			av_debugaccess        => open,                                                                              --              (terminated)
			av_outputenable       => open                                                                               --              (terminated)
		);

	no_of_cam_channels_s1_translator : component de4_qsys_button_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => clk_clk,                                                                          --                      clk.clk
			reset                 => rst_controller_001_reset_out_reset,                                               --                    reset.reset
			uav_address           => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => no_of_cam_channels_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => no_of_cam_channels_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => no_of_cam_channels_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => no_of_cam_channels_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => no_of_cam_channels_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read               => open,                                                                             --              (terminated)
			av_begintransfer      => open,                                                                             --              (terminated)
			av_beginbursttransfer => open,                                                                             --              (terminated)
			av_burstcount         => open,                                                                             --              (terminated)
			av_byteenable         => open,                                                                             --              (terminated)
			av_readdatavalid      => '0',                                                                              --              (terminated)
			av_waitrequest        => '0',                                                                              --              (terminated)
			av_writebyteenable    => open,                                                                             --              (terminated)
			av_lock               => open,                                                                             --              (terminated)
			av_clken              => open,                                                                             --              (terminated)
			uav_clken             => '0',                                                                              --              (terminated)
			av_debugaccess        => open,                                                                             --              (terminated)
			av_outputenable       => open                                                                              --              (terminated)
		);

	nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent : component DE4_QSYS_nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => mem_if_ddr2_emif_afi_clk_clk,                                                              --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			av_address       => nios2_qsys_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => limiter_rsp_src_valid,                                                                     --        rp.valid
			rp_data          => limiter_rsp_src_data,                                                                      --          .data
			rp_channel       => limiter_rsp_src_channel,                                                                   --          .channel
			rp_startofpacket => limiter_rsp_src_startofpacket,                                                             --          .startofpacket
			rp_endofpacket   => limiter_rsp_src_endofpacket,                                                               --          .endofpacket
			rp_ready         => limiter_rsp_src_ready                                                                      --          .ready
		);

	nios2_qsys_data_master_translator_avalon_universal_master_0_agent : component DE4_QSYS_nios2_qsys_data_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => mem_if_ddr2_emif_afi_clk_clk,                                                       --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address       => nios2_qsys_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => nios2_qsys_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => nios2_qsys_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => nios2_qsys_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => nios2_qsys_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => nios2_qsys_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => limiter_001_rsp_src_valid,                                                          --        rp.valid
			rp_data          => limiter_001_rsp_src_data,                                                           --          .data
			rp_channel       => limiter_001_rsp_src_channel,                                                        --          .channel
			rp_startofpacket => limiter_001_rsp_src_startofpacket,                                                  --          .startofpacket
			rp_endofpacket   => limiter_001_rsp_src_endofpacket,                                                    --          .endofpacket
			rp_ready         => limiter_001_rsp_src_ready                                                           --          .ready
		);

	mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent : component DE4_QSYS_mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent
		port map (
			clk              => mem_if_ddr2_emif_afi_clk_clk,                                                               --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			av_address       => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => limiter_002_rsp_src_valid,                                                                  --        rp.valid
			rp_data          => limiter_002_rsp_src_data,                                                                   --          .data
			rp_channel       => limiter_002_rsp_src_channel,                                                                --          .channel
			rp_startofpacket => limiter_002_rsp_src_startofpacket,                                                          --          .startofpacket
			rp_endofpacket   => limiter_002_rsp_src_endofpacket,                                                            --          .endofpacket
			rp_ready         => limiter_002_rsp_src_ready                                                                   --          .ready
		);

	dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent : component DE4_QSYS_dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => mem_if_ddr2_emif_afi_clk_clk,                                                                     --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			av_address       => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => width_adapter_004_src_valid,                                                                      --        rp.valid
			rp_data          => width_adapter_004_src_data,                                                                       --          .data
			rp_channel       => width_adapter_004_src_channel,                                                                    --          .channel
			rp_startofpacket => width_adapter_004_src_startofpacket,                                                              --          .startofpacket
			rp_endofpacket   => width_adapter_004_src_endofpacket,                                                                --          .endofpacket
			rp_ready         => width_adapter_004_src_ready                                                                       --          .ready
		);

	cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent : component DE4_QSYS_cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => mem_if_ddr2_emif_afi_clk_clk,                                                                     --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			av_address       => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => width_adapter_005_src_valid,                                                                      --        rp.valid
			rp_data          => width_adapter_005_src_data,                                                                       --          .data
			rp_channel       => width_adapter_005_src_channel,                                                                    --          .channel
			rp_startofpacket => width_adapter_005_src_startofpacket,                                                              --          .startofpacket
			rp_endofpacket   => width_adapter_005_src_endofpacket,                                                                --          .endofpacket
			rp_ready         => width_adapter_005_src_ready                                                                       --          .ready
		);

	nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => mem_if_ddr2_emif_afi_clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                    --       clk_reset.reset
			m0_address              => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                       --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                       --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                        --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                                 --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                                     --                .channel
			rf_sink_ready           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                    -- clk_reset.reset
			in_data           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent : component DE4_QSYS_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => mem_if_ddr2_emif_afi_clk_clk,                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                       --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                       --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                        --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                                 --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                     --                .channel
			rf_sink_ready           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component DE4_QSYS_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => mem_if_ddr2_emif_afi_clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_002_source0_ready,                                                                  --              cp.ready
			cp_valid                => burst_adapter_002_source0_valid,                                                                  --                .valid
			cp_data                 => burst_adapter_002_source0_data,                                                                   --                .data
			cp_startofpacket        => burst_adapter_002_source0_startofpacket,                                                          --                .startofpacket
			cp_endofpacket          => burst_adapter_002_source0_endofpacket,                                                            --                .endofpacket
			cp_channel              => burst_adapter_002_source0_channel,                                                                --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent : component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                             --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                  --       clk_reset.reset
			m0_address              => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_003_source0_ready,                                                                     --              cp.ready
			cp_valid                => burst_adapter_003_source0_valid,                                                                     --                .valid
			cp_data                 => burst_adapter_003_source0_data,                                                                      --                .data
			cp_startofpacket        => burst_adapter_003_source0_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => burst_adapter_003_source0_endofpacket,                                                               --                .endofpacket
			cp_channel              => burst_adapter_003_source0_channel,                                                                   --                .channel
			rf_sink_ready           => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                             --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                  -- clk_reset.reset
			in_data           => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                                       --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                                            -- clk_reset.reset
			in_data   => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	button_s1_translator_avalon_universal_slave_0_agent : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                        --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                             --       clk_reset.reset
			m0_address              => button_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => button_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => button_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => button_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => button_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => button_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => button_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => button_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => button_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_004_source0_ready,                                                --              cp.ready
			cp_valid                => burst_adapter_004_source0_valid,                                                --                .valid
			cp_data                 => burst_adapter_004_source0_data,                                                 --                .data
			cp_startofpacket        => burst_adapter_004_source0_startofpacket,                                        --                .startofpacket
			cp_endofpacket          => burst_adapter_004_source0_endofpacket,                                          --                .endofpacket
			cp_channel              => burst_adapter_004_source0_channel,                                              --                .channel
			rf_sink_ready           => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => button_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                        --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			in_data           => button_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                  --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                       -- clk_reset.reset
			in_data   => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	led_s1_translator_avalon_universal_slave_0_agent : component DE4_QSYS_led_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                          --       clk_reset.reset
			m0_address              => led_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => led_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => led_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => led_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => led_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => led_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => led_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => led_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => led_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_005_source0_ready,                                             --              cp.ready
			cp_valid                => burst_adapter_005_source0_valid,                                             --                .valid
			cp_data                 => burst_adapter_005_source0_data,                                              --                .data
			cp_startofpacket        => burst_adapter_005_source0_startofpacket,                                     --                .startofpacket
			cp_endofpacket          => burst_adapter_005_source0_endofpacket,                                       --                .endofpacket
			cp_channel              => burst_adapter_005_source0_channel,                                           --                .channel
			rf_sink_ready           => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			in_data           => led_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                               --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                    -- clk_reset.reset
			in_data   => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	timer_s1_translator_avalon_universal_slave_0_agent : component DE4_QSYS_timer_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                       --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                            --       clk_reset.reset
			m0_address              => timer_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_006_source0_ready,                                               --              cp.ready
			cp_valid                => burst_adapter_006_source0_valid,                                               --                .valid
			cp_data                 => burst_adapter_006_source0_data,                                                --                .data
			cp_startofpacket        => burst_adapter_006_source0_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => burst_adapter_006_source0_endofpacket,                                         --                .endofpacket
			cp_channel              => burst_adapter_006_source0_channel,                                             --                .channel
			rf_sink_ready           => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                       --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			in_data           => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                 --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                      -- clk_reset.reset
			in_data   => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	spi_2_spi_control_port_translator_avalon_universal_slave_0_agent : component DE4_QSYS_spi_2_spi_control_port_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_007_source0_ready,                                                             --              cp.ready
			cp_valid                => burst_adapter_007_source0_valid,                                                             --                .valid
			cp_data                 => burst_adapter_007_source0_data,                                                              --                .data
			cp_startofpacket        => burst_adapter_007_source0_startofpacket,                                                     --                .startofpacket
			cp_endofpacket          => burst_adapter_007_source0_endofpacket,                                                       --                .endofpacket
			cp_channel              => burst_adapter_007_source0_channel,                                                           --                .channel
			rf_sink_ready           => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                               --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                                    -- clk_reset.reset
			in_data   => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component DE4_QSYS_sysid_control_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                       --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_008_source0_ready,                                                          --              cp.ready
			cp_valid                => burst_adapter_008_source0_valid,                                                          --                .valid
			cp_data                 => burst_adapter_008_source0_data,                                                           --                .data
			cp_startofpacket        => burst_adapter_008_source0_startofpacket,                                                  --                .startofpacket
			cp_endofpacket          => burst_adapter_008_source0_endofpacket,                                                    --                .endofpacket
			cp_channel              => burst_adapter_008_source0_channel,                                                        --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                            --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			in_data   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent : component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => mem_if_ddr2_emif_afi_clk_clk,                                                              --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_009_src_ready,                                                                --              cp.ready
			cp_valid                => cmd_xbar_mux_009_src_valid,                                                                --                .valid
			cp_data                 => cmd_xbar_mux_009_src_data,                                                                 --                .data
			cp_startofpacket        => cmd_xbar_mux_009_src_startofpacket,                                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_009_src_endofpacket,                                                          --                .endofpacket
			cp_channel              => cmd_xbar_mux_009_src_channel,                                                              --                .channel
			rf_sink_ready           => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,                                                              --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => mem_if_ddr2_emif_afi_clk_clk,                                                        --       clk.clk
			reset     => rst_controller_002_reset_out_reset,                                                  -- clk_reset.reset
			in_data   => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	spi_1_spi_control_port_translator_avalon_universal_slave_0_agent : component DE4_QSYS_spi_1_spi_control_port_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_009_source0_ready,                                                             --              cp.ready
			cp_valid                => burst_adapter_009_source0_valid,                                                             --                .valid
			cp_data                 => burst_adapter_009_source0_data,                                                              --                .data
			cp_startofpacket        => burst_adapter_009_source0_startofpacket,                                                     --                .startofpacket
			cp_endofpacket          => burst_adapter_009_source0_endofpacket,                                                       --                .endofpacket
			cp_channel              => burst_adapter_009_source0_channel,                                                           --                .channel
			rf_sink_ready           => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                               --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                                    -- clk_reset.reset
			in_data   => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent : component DE4_QSYS_no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                    --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_010_source0_ready,                                                            --              cp.ready
			cp_valid                => burst_adapter_010_source0_valid,                                                            --                .valid
			cp_data                 => burst_adapter_010_source0_data,                                                             --                .data
			cp_startofpacket        => burst_adapter_010_source0_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => burst_adapter_010_source0_endofpacket,                                                      --                .endofpacket
			cp_channel              => burst_adapter_010_source0_channel,                                                          --                .channel
			rf_sink_ready           => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component DE4_QSYS_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component DE4_QSYS_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                              --       clk.clk
			reset     => rst_controller_001_reset_out_reset,                                                   -- clk_reset.reset
			in_data   => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	addr_router : component DE4_QSYS_addr_router
		port map (
			sink_ready         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                     --       src.ready
			src_valid          => addr_router_src_valid,                                                                     --          .valid
			src_data           => addr_router_src_data,                                                                      --          .data
			src_channel        => addr_router_src_channel,                                                                   --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                --          .endofpacket
		);

	addr_router_001 : component DE4_QSYS_addr_router_001
		port map (
			sink_ready         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                       --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                          --       src.ready
			src_valid          => addr_router_001_src_valid,                                                          --          .valid
			src_data           => addr_router_001_src_data,                                                           --          .data
			src_channel        => addr_router_001_src_channel,                                                        --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                     --          .endofpacket
		);

	addr_router_002 : component DE4_QSYS_addr_router_002
		port map (
			sink_ready         => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			src_ready          => addr_router_002_src_ready,                                                                  --       src.ready
			src_valid          => addr_router_002_src_valid,                                                                  --          .valid
			src_data           => addr_router_002_src_data,                                                                   --          .data
			src_channel        => addr_router_002_src_channel,                                                                --          .channel
			src_startofpacket  => addr_router_002_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => addr_router_002_src_endofpacket                                                             --          .endofpacket
		);

	addr_router_003 : component DE4_QSYS_addr_router_003
		port map (
			sink_ready         => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => dvi_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			src_ready          => addr_router_003_src_ready,                                                                        --       src.ready
			src_valid          => addr_router_003_src_valid,                                                                        --          .valid
			src_data           => addr_router_003_src_data,                                                                         --          .data
			src_channel        => addr_router_003_src_channel,                                                                      --          .channel
			src_startofpacket  => addr_router_003_src_startofpacket,                                                                --          .startofpacket
			src_endofpacket    => addr_router_003_src_endofpacket                                                                   --          .endofpacket
		);

	addr_router_004 : component DE4_QSYS_addr_router_004
		port map (
			sink_ready         => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cmv_master_interface_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			src_ready          => addr_router_004_src_ready,                                                                        --       src.ready
			src_valid          => addr_router_004_src_valid,                                                                        --          .valid
			src_data           => addr_router_004_src_data,                                                                         --          .data
			src_channel        => addr_router_004_src_channel,                                                                      --          .channel
			src_startofpacket  => addr_router_004_src_startofpacket,                                                                --          .startofpacket
			src_endofpacket    => addr_router_004_src_endofpacket                                                                   --          .endofpacket
		);

	id_router : component DE4_QSYS_id_router
		port map (
			sink_ready         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                     --       src.ready
			src_valid          => id_router_src_valid,                                                                     --          .valid
			src_data           => id_router_src_data,                                                                      --          .data
			src_channel        => id_router_src_channel,                                                                   --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                                --          .endofpacket
		);

	id_router_001 : component DE4_QSYS_id_router
		port map (
			sink_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                     --       src.ready
			src_valid          => id_router_001_src_valid,                                                     --          .valid
			src_data           => id_router_001_src_data,                                                      --          .data
			src_channel        => id_router_001_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                --          .endofpacket
		);

	id_router_002 : component DE4_QSYS_id_router_002
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                --       src.ready
			src_valid          => id_router_002_src_valid,                                                                --          .valid
			src_data           => id_router_002_src_data,                                                                 --          .data
			src_channel        => id_router_002_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                           --          .endofpacket
		);

	id_router_003 : component DE4_QSYS_id_router_002
		port map (
			sink_ready         => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                                   --       src.ready
			src_valid          => id_router_003_src_valid,                                                                   --          .valid
			src_data           => id_router_003_src_data,                                                                    --          .data
			src_channel        => id_router_003_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                              --          .endofpacket
		);

	id_router_004 : component DE4_QSYS_id_router_004
		port map (
			sink_ready         => button_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => button_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => button_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                              --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                   -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                              --       src.ready
			src_valid          => id_router_004_src_valid,                                              --          .valid
			src_data           => id_router_004_src_data,                                               --          .data
			src_channel        => id_router_004_src_channel,                                            --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                         --          .endofpacket
		);

	id_router_005 : component DE4_QSYS_id_router_004
		port map (
			sink_ready         => led_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => led_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => led_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                           --       src.ready
			src_valid          => id_router_005_src_valid,                                           --          .valid
			src_data           => id_router_005_src_data,                                            --          .data
			src_channel        => id_router_005_src_channel,                                         --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                      --          .endofpacket
		);

	id_router_006 : component DE4_QSYS_id_router_004
		port map (
			sink_ready         => timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                             --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                  -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                             --       src.ready
			src_valid          => id_router_006_src_valid,                                             --          .valid
			src_data           => id_router_006_src_data,                                              --          .data
			src_channel        => id_router_006_src_channel,                                           --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                        --          .endofpacket
		);

	id_router_007 : component DE4_QSYS_id_router_004
		port map (
			sink_ready         => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => spi_2_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                           --       src.ready
			src_valid          => id_router_007_src_valid,                                                           --          .valid
			src_data           => id_router_007_src_data,                                                            --          .data
			src_channel        => id_router_007_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                      --          .endofpacket
		);

	id_router_008 : component DE4_QSYS_id_router_004
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                        --       src.ready
			src_valid          => id_router_008_src_valid,                                                        --          .valid
			src_data           => id_router_008_src_data,                                                         --          .data
			src_channel        => id_router_008_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                   --          .endofpacket
		);

	id_router_009 : component DE4_QSYS_id_router_009
		port map (
			sink_ready         => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => mem_if_ddr2_emif_afi_clk_clk,                                                    --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                         --       src.ready
			src_valid          => id_router_009_src_valid,                                                         --          .valid
			src_data           => id_router_009_src_data,                                                          --          .data
			src_channel        => id_router_009_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                    --          .endofpacket
		);

	id_router_010 : component DE4_QSYS_id_router_004
		port map (
			sink_ready         => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => spi_1_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                                           --       src.ready
			src_valid          => id_router_010_src_valid,                                                           --          .valid
			src_data           => id_router_010_src_data,                                                            --          .data
			src_channel        => id_router_010_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                                      --          .endofpacket
		);

	id_router_011 : component DE4_QSYS_id_router_004
		port map (
			sink_ready         => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => no_of_cam_channels_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                          --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                          --       src.ready
			src_valid          => id_router_011_src_valid,                                                          --          .valid
			src_data           => id_router_011_src_data,                                                           --          .data
			src_channel        => id_router_011_src_channel,                                                        --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                                     --          .endofpacket
		);

	limiter : component DE4_QSYS_limiter
		port map (
			clk                    => mem_if_ddr2_emif_afi_clk_clk,   --       clk.clk
			reset                  => rst_controller_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,          --          .valid
			cmd_sink_data          => addr_router_src_data,           --          .data
			cmd_sink_channel       => addr_router_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data          -- cmd_valid.data
		);

	limiter_001 : component DE4_QSYS_limiter_001
		port map (
			clk                    => mem_if_ddr2_emif_afi_clk_clk,       --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_001_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_001_src_valid,          --          .valid
			cmd_sink_data          => addr_router_001_src_data,           --          .data
			cmd_sink_channel       => addr_router_001_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_001_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_001_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_001_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_001_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_001_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_001_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_001_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_001_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_001_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_001_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_001_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_001_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_001_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_001_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_001_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_001_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_001_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_001_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_001_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_001_cmd_valid_data          -- cmd_valid.data
		);

	limiter_002 : component DE4_QSYS_limiter_002
		port map (
			clk                    => mem_if_ddr2_emif_afi_clk_clk,       --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_002_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_002_src_valid,          --          .valid
			cmd_sink_data          => addr_router_002_src_data,           --          .data
			cmd_sink_channel       => addr_router_002_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_002_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_002_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_002_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_002_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_002_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_002_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_002_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_002_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_002_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_002_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_002_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_002_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_002_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_002_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_002_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_002_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_002_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_002_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_002_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_002_cmd_valid_data          -- cmd_valid.data
		);

	burst_adapter : component DE4_QSYS_burst_adapter
		port map (
			clk                   => mem_if_ddr2_emif_afi_clk_clk,        --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_src_ready,              --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component DE4_QSYS_burst_adapter
		port map (
			clk                   => mem_if_ddr2_emif_afi_clk_clk,            --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_001_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_001_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_001_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_001_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_001_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_001_src_ready,              --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	burst_adapter_002 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => mem_if_ddr2_emif_afi_clk_clk,            --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => cmd_xbar_demux_001_src2_valid,           --     sink0.valid
			sink0_data            => cmd_xbar_demux_001_src2_data,            --          .data
			sink0_channel         => cmd_xbar_demux_001_src2_channel,         --          .channel
			sink0_startofpacket   => cmd_xbar_demux_001_src2_startofpacket,   --          .startofpacket
			sink0_endofpacket     => cmd_xbar_demux_001_src2_endofpacket,     --          .endofpacket
			sink0_ready           => cmd_xbar_demux_001_src2_ready,           --          .ready
			source0_valid         => burst_adapter_002_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_002_source0_data,          --          .data
			source0_channel       => burst_adapter_002_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_002_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_002_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_002_source0_ready          --          .ready
		);

	burst_adapter_003 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => crosser_out_valid,                       --     sink0.valid
			sink0_data            => crosser_out_data,                        --          .data
			sink0_channel         => crosser_out_channel,                     --          .channel
			sink0_startofpacket   => crosser_out_startofpacket,               --          .startofpacket
			sink0_endofpacket     => crosser_out_endofpacket,                 --          .endofpacket
			sink0_ready           => crosser_out_ready,                       --          .ready
			source0_valid         => burst_adapter_003_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_003_source0_data,          --          .data
			source0_channel       => burst_adapter_003_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_003_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_003_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_003_source0_ready          --          .ready
		);

	burst_adapter_004 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_004_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_004_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_004_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_004_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_004_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_004_src_ready,              --          .ready
			source0_valid         => burst_adapter_004_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_004_source0_data,          --          .data
			source0_channel       => burst_adapter_004_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_004_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_004_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_004_source0_ready          --          .ready
		);

	burst_adapter_005 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_005_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_005_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_005_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_005_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_005_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_005_src_ready,              --          .ready
			source0_valid         => burst_adapter_005_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_005_source0_data,          --          .data
			source0_channel       => burst_adapter_005_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_005_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_005_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_005_source0_ready          --          .ready
		);

	burst_adapter_006 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_006_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_006_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_006_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_006_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_006_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_006_src_ready,              --          .ready
			source0_valid         => burst_adapter_006_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_006_source0_data,          --          .data
			source0_channel       => burst_adapter_006_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_006_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_006_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_006_source0_ready          --          .ready
		);

	burst_adapter_007 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_007_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_007_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_007_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_007_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_007_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_007_src_ready,              --          .ready
			source0_valid         => burst_adapter_007_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_007_source0_data,          --          .data
			source0_channel       => burst_adapter_007_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_007_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_007_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_007_source0_ready          --          .ready
		);

	burst_adapter_008 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_008_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_008_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_008_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_008_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_008_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_008_src_ready,              --          .ready
			source0_valid         => burst_adapter_008_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_008_source0_data,          --          .data
			source0_channel       => burst_adapter_008_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_008_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_008_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_008_source0_ready          --          .ready
		);

	burst_adapter_009 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_010_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_010_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_010_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_010_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_010_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_010_src_ready,              --          .ready
			source0_valid         => burst_adapter_009_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_009_source0_data,          --          .data
			source0_channel       => burst_adapter_009_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_009_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_009_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_009_source0_ready          --          .ready
		);

	burst_adapter_010 : component DE4_QSYS_burst_adapter_002
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_011_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_011_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_011_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_011_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_011_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_011_src_ready,              --          .ready
			source0_valid         => burst_adapter_010_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_010_source0_data,          --          .data
			source0_channel       => burst_adapter_010_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_010_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_010_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_010_source0_ready          --          .ready
		);

	rst_controller : component DE4_QSYS_rst_controller
		port map (
			reset_in0 => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk       => mem_if_ddr2_emif_afi_clk_clk,   --       clk.clk
			reset_out => rst_controller_reset_out_reset  -- reset_out.reset
		);

	rst_controller_001 : component DE4_QSYS_rst_controller
		port map (
			reset_in0 => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk       => clk_clk,                            --       clk.clk
			reset_out => rst_controller_001_reset_out_reset  -- reset_out.reset
		);

	rst_controller_002 : component DE4_QSYS_rst_controller
		port map (
			reset_in0 => mem_if_ddr2_emif_afi_reset_reset_ports_inv, -- reset_in0.reset
			clk       => mem_if_ddr2_emif_afi_clk_clk,               --       clk.clk
			reset_out => rst_controller_002_reset_out_reset          -- reset_out.reset
		);

	cmd_xbar_demux : component DE4_QSYS_cmd_xbar_demux
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,      --        clk.clk
			reset              => rst_controller_reset_out_reset,    --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_cmd_src_channel,           --           .channel
			sink_data          => limiter_cmd_src_data,              --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_001 : component DE4_QSYS_cmd_xbar_demux_001
		port map (
			clk                 => mem_if_ddr2_emif_afi_clk_clk,           --        clk.clk
			reset               => rst_controller_reset_out_reset,         --  clk_reset.reset
			sink_ready          => limiter_001_cmd_src_ready,              --       sink.ready
			sink_channel        => limiter_001_cmd_src_channel,            --           .channel
			sink_data           => limiter_001_cmd_src_data,               --           .data
			sink_startofpacket  => limiter_001_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket    => limiter_001_cmd_src_endofpacket,        --           .endofpacket
			sink_valid          => limiter_001_cmd_valid_data,             -- sink_valid.data
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --       src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --           .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --           .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --           .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --           .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --           .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --       src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --           .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --           .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --           .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --           .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --           .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --       src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --           .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --           .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --           .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --           .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --           .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --       src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --           .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --           .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --           .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --           .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --           .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --       src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --           .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --           .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --           .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --           .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --           .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --       src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --           .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --           .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --           .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --           .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --           .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --       src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --           .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --           .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --           .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --           .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --           .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --       src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --           .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --           .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --           .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --           .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --           .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --       src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --           .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --           .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --           .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --           .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --           .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --       src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --           .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --           .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --           .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --           .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --           .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --      src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --           .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --           .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --           .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --           .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket,   --           .endofpacket
			src11_ready         => cmd_xbar_demux_001_src11_ready,         --      src11.ready
			src11_valid         => cmd_xbar_demux_001_src11_valid,         --           .valid
			src11_data          => cmd_xbar_demux_001_src11_data,          --           .data
			src11_channel       => cmd_xbar_demux_001_src11_channel,       --           .channel
			src11_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --           .startofpacket
			src11_endofpacket   => cmd_xbar_demux_001_src11_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_002 : component DE4_QSYS_cmd_xbar_demux_002
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,          --        clk.clk
			reset              => rst_controller_reset_out_reset,        --  clk_reset.reset
			sink_ready         => limiter_002_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_002_cmd_src_channel,           --           .channel
			sink_data          => limiter_002_cmd_src_data,              --           .data
			sink_startofpacket => limiter_002_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_002_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_002_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_002_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_002_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_002_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_002_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_002_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_002_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_002_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_002_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_002_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_002_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_002_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_002_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_002_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_002_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_002_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_002_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_002_src2_endofpacket,   --           .endofpacket
			src3_ready         => cmd_xbar_demux_002_src3_ready,         --       src3.ready
			src3_valid         => cmd_xbar_demux_002_src3_valid,         --           .valid
			src3_data          => cmd_xbar_demux_002_src3_data,          --           .data
			src3_channel       => cmd_xbar_demux_002_src3_channel,       --           .channel
			src3_startofpacket => cmd_xbar_demux_002_src3_startofpacket, --           .startofpacket
			src3_endofpacket   => cmd_xbar_demux_002_src3_endofpacket,   --           .endofpacket
			src4_ready         => cmd_xbar_demux_002_src4_ready,         --       src4.ready
			src4_valid         => cmd_xbar_demux_002_src4_valid,         --           .valid
			src4_data          => cmd_xbar_demux_002_src4_data,          --           .data
			src4_channel       => cmd_xbar_demux_002_src4_channel,       --           .channel
			src4_startofpacket => cmd_xbar_demux_002_src4_startofpacket, --           .startofpacket
			src4_endofpacket   => cmd_xbar_demux_002_src4_endofpacket,   --           .endofpacket
			src5_ready         => cmd_xbar_demux_002_src5_ready,         --       src5.ready
			src5_valid         => cmd_xbar_demux_002_src5_valid,         --           .valid
			src5_data          => cmd_xbar_demux_002_src5_data,          --           .data
			src5_channel       => cmd_xbar_demux_002_src5_channel,       --           .channel
			src5_startofpacket => cmd_xbar_demux_002_src5_startofpacket, --           .startofpacket
			src5_endofpacket   => cmd_xbar_demux_002_src5_endofpacket,   --           .endofpacket
			src6_ready         => cmd_xbar_demux_002_src6_ready,         --       src6.ready
			src6_valid         => cmd_xbar_demux_002_src6_valid,         --           .valid
			src6_data          => cmd_xbar_demux_002_src6_data,          --           .data
			src6_channel       => cmd_xbar_demux_002_src6_channel,       --           .channel
			src6_startofpacket => cmd_xbar_demux_002_src6_startofpacket, --           .startofpacket
			src6_endofpacket   => cmd_xbar_demux_002_src6_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_003 : component DE4_QSYS_cmd_xbar_demux_003
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_003_src_ready,             --      sink.ready
			sink_channel       => addr_router_003_src_channel,           --          .channel
			sink_data          => addr_router_003_src_data,              --          .data
			sink_startofpacket => addr_router_003_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_003_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_003_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_003_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_004 : component DE4_QSYS_cmd_xbar_demux_004
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_004_src_ready,             --      sink.ready
			sink_channel       => addr_router_004_src_channel,           --          .channel
			sink_data          => addr_router_004_src_data,              --          .data
			sink_startofpacket => addr_router_004_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_004_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_004_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_004_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_001_reset_out_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,         --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,         --          .valid
			src_data            => cmd_xbar_mux_004_src_data,          --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,       --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket, --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_001_out_ready,              --     sink0.ready
			sink0_valid         => crosser_001_out_valid,              --          .valid
			sink0_channel       => crosser_001_out_channel,            --          .channel
			sink0_data          => crosser_001_out_data,               --          .data
			sink0_startofpacket => crosser_001_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_001_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_008_out_ready,              --     sink1.ready
			sink1_valid         => crosser_008_out_valid,              --          .valid
			sink1_channel       => crosser_008_out_channel,            --          .channel
			sink1_data          => crosser_008_out_data,               --          .data
			sink1_startofpacket => crosser_008_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_008_out_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_005 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_001_reset_out_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_005_src_ready,         --       src.ready
			src_valid           => cmd_xbar_mux_005_src_valid,         --          .valid
			src_data            => cmd_xbar_mux_005_src_data,          --          .data
			src_channel         => cmd_xbar_mux_005_src_channel,       --          .channel
			src_startofpacket   => cmd_xbar_mux_005_src_startofpacket, --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_005_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_002_out_ready,              --     sink0.ready
			sink0_valid         => crosser_002_out_valid,              --          .valid
			sink0_channel       => crosser_002_out_channel,            --          .channel
			sink0_data          => crosser_002_out_data,               --          .data
			sink0_startofpacket => crosser_002_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_002_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_009_out_ready,              --     sink1.ready
			sink1_valid         => crosser_009_out_valid,              --          .valid
			sink1_channel       => crosser_009_out_channel,            --          .channel
			sink1_data          => crosser_009_out_data,               --          .data
			sink1_startofpacket => crosser_009_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_009_out_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_006 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_001_reset_out_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_006_src_ready,         --       src.ready
			src_valid           => cmd_xbar_mux_006_src_valid,         --          .valid
			src_data            => cmd_xbar_mux_006_src_data,          --          .data
			src_channel         => cmd_xbar_mux_006_src_channel,       --          .channel
			src_startofpacket   => cmd_xbar_mux_006_src_startofpacket, --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_006_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_003_out_ready,              --     sink0.ready
			sink0_valid         => crosser_003_out_valid,              --          .valid
			sink0_channel       => crosser_003_out_channel,            --          .channel
			sink0_data          => crosser_003_out_data,               --          .data
			sink0_startofpacket => crosser_003_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_003_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_010_out_ready,              --     sink1.ready
			sink1_valid         => crosser_010_out_valid,              --          .valid
			sink1_channel       => crosser_010_out_channel,            --          .channel
			sink1_data          => crosser_010_out_data,               --          .data
			sink1_startofpacket => crosser_010_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_010_out_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_007 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_001_reset_out_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_007_src_ready,         --       src.ready
			src_valid           => cmd_xbar_mux_007_src_valid,         --          .valid
			src_data            => cmd_xbar_mux_007_src_data,          --          .data
			src_channel         => cmd_xbar_mux_007_src_channel,       --          .channel
			src_startofpacket   => cmd_xbar_mux_007_src_startofpacket, --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_007_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_004_out_ready,              --     sink0.ready
			sink0_valid         => crosser_004_out_valid,              --          .valid
			sink0_channel       => crosser_004_out_channel,            --          .channel
			sink0_data          => crosser_004_out_data,               --          .data
			sink0_startofpacket => crosser_004_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_004_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_011_out_ready,              --     sink1.ready
			sink1_valid         => crosser_011_out_valid,              --          .valid
			sink1_channel       => crosser_011_out_channel,            --          .channel
			sink1_data          => crosser_011_out_data,               --          .data
			sink1_startofpacket => crosser_011_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_011_out_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_008 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_001_reset_out_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_008_src_ready,         --       src.ready
			src_valid           => cmd_xbar_mux_008_src_valid,         --          .valid
			src_data            => cmd_xbar_mux_008_src_data,          --          .data
			src_channel         => cmd_xbar_mux_008_src_channel,       --          .channel
			src_startofpacket   => cmd_xbar_mux_008_src_startofpacket, --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_008_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_005_out_ready,              --     sink0.ready
			sink0_valid         => crosser_005_out_valid,              --          .valid
			sink0_channel       => crosser_005_out_channel,            --          .channel
			sink0_data          => crosser_005_out_data,               --          .data
			sink0_startofpacket => crosser_005_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_005_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_012_out_ready,              --     sink1.ready
			sink1_valid         => crosser_012_out_valid,              --          .valid
			sink1_channel       => crosser_012_out_channel,            --          .channel
			sink1_data          => crosser_012_out_data,               --          .data
			sink1_startofpacket => crosser_012_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_012_out_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_009 : component DE4_QSYS_cmd_xbar_mux_009
		port map (
			clk                 => mem_if_ddr2_emif_afi_clk_clk,        --       clk.clk
			reset               => rst_controller_002_reset_out_reset,  -- clk_reset.reset
			src_ready           => cmd_xbar_mux_009_src_ready,          --       src.ready
			src_valid           => cmd_xbar_mux_009_src_valid,          --          .valid
			src_data            => cmd_xbar_mux_009_src_data,           --          .data
			src_channel         => cmd_xbar_mux_009_src_channel,        --          .channel
			src_startofpacket   => cmd_xbar_mux_009_src_startofpacket,  --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_009_src_endofpacket,    --          .endofpacket
			sink0_ready         => width_adapter_src_ready,             --     sink0.ready
			sink0_valid         => width_adapter_src_valid,             --          .valid
			sink0_channel       => width_adapter_src_channel,           --          .channel
			sink0_data          => width_adapter_src_data,              --          .data
			sink0_startofpacket => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket   => width_adapter_src_endofpacket,       --          .endofpacket
			sink1_ready         => width_adapter_001_src_ready,         --     sink1.ready
			sink1_valid         => width_adapter_001_src_valid,         --          .valid
			sink1_channel       => width_adapter_001_src_channel,       --          .channel
			sink1_data          => width_adapter_001_src_data,          --          .data
			sink1_startofpacket => width_adapter_001_src_startofpacket, --          .startofpacket
			sink1_endofpacket   => width_adapter_001_src_endofpacket,   --          .endofpacket
			sink2_ready         => width_adapter_002_src_ready,         --     sink2.ready
			sink2_valid         => width_adapter_002_src_valid,         --          .valid
			sink2_channel       => width_adapter_002_src_channel,       --          .channel
			sink2_data          => width_adapter_002_src_data,          --          .data
			sink2_startofpacket => width_adapter_002_src_startofpacket, --          .startofpacket
			sink2_endofpacket   => width_adapter_002_src_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_010 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_001_reset_out_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_010_src_ready,         --       src.ready
			src_valid           => cmd_xbar_mux_010_src_valid,         --          .valid
			src_data            => cmd_xbar_mux_010_src_data,          --          .data
			src_channel         => cmd_xbar_mux_010_src_channel,       --          .channel
			src_startofpacket   => cmd_xbar_mux_010_src_startofpacket, --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_010_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_006_out_ready,              --     sink0.ready
			sink0_valid         => crosser_006_out_valid,              --          .valid
			sink0_channel       => crosser_006_out_channel,            --          .channel
			sink0_data          => crosser_006_out_data,               --          .data
			sink0_startofpacket => crosser_006_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_006_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_013_out_ready,              --     sink1.ready
			sink1_valid         => crosser_013_out_valid,              --          .valid
			sink1_channel       => crosser_013_out_channel,            --          .channel
			sink1_data          => crosser_013_out_data,               --          .data
			sink1_startofpacket => crosser_013_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_013_out_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_011 : component DE4_QSYS_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_001_reset_out_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_011_src_ready,         --       src.ready
			src_valid           => cmd_xbar_mux_011_src_valid,         --          .valid
			src_data            => cmd_xbar_mux_011_src_data,          --          .data
			src_channel         => cmd_xbar_mux_011_src_channel,       --          .channel
			src_startofpacket   => cmd_xbar_mux_011_src_startofpacket, --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_011_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_007_out_ready,              --     sink0.ready
			sink0_valid         => crosser_007_out_valid,              --          .valid
			sink0_channel       => crosser_007_out_channel,            --          .channel
			sink0_data          => crosser_007_out_data,               --          .data
			sink0_startofpacket => crosser_007_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_007_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_014_out_ready,              --     sink1.ready
			sink1_valid         => crosser_014_out_valid,              --          .valid
			sink1_channel       => crosser_014_out_channel,            --          .channel
			sink1_data          => crosser_014_out_data,               --          .data
			sink1_startofpacket => crosser_014_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_014_out_endofpacket         --          .endofpacket
		);

	rsp_xbar_demux : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,      --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component DE4_QSYS_cmd_xbar_demux_003
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component DE4_QSYS_cmd_xbar_demux_003
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_005_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_005_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_005_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_005_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_005_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_006_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_006_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_006_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_006_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_006_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_007_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_007_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_007_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_007_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_007_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_007_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_008_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_008_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_008_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_008_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_008_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_008_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component DE4_QSYS_rsp_xbar_demux_009
		port map (
			clk                => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_009_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_009_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_009_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_009_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_009_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_009_src1_endofpacket,   --          .endofpacket
			src2_ready         => rsp_xbar_demux_009_src2_ready,         --      src2.ready
			src2_valid         => rsp_xbar_demux_009_src2_valid,         --          .valid
			src2_data          => rsp_xbar_demux_009_src2_data,          --          .data
			src2_channel       => rsp_xbar_demux_009_src2_channel,       --          .channel
			src2_startofpacket => rsp_xbar_demux_009_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => rsp_xbar_demux_009_src2_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_010_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_010_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_010_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_010_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_010_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_010_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component DE4_QSYS_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_011_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_011_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_011_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_011_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_011_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_011_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component DE4_QSYS_rsp_xbar_mux
		port map (
			clk                 => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component DE4_QSYS_rsp_xbar_mux_001
		port map (
			clk                  => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready          => crosser_015_out_ready,                 --     sink3.ready
			sink3_valid          => crosser_015_out_valid,                 --          .valid
			sink3_channel        => crosser_015_out_channel,               --          .channel
			sink3_data           => crosser_015_out_data,                  --          .data
			sink3_startofpacket  => crosser_015_out_startofpacket,         --          .startofpacket
			sink3_endofpacket    => crosser_015_out_endofpacket,           --          .endofpacket
			sink4_ready          => crosser_016_out_ready,                 --     sink4.ready
			sink4_valid          => crosser_016_out_valid,                 --          .valid
			sink4_channel        => crosser_016_out_channel,               --          .channel
			sink4_data           => crosser_016_out_data,                  --          .data
			sink4_startofpacket  => crosser_016_out_startofpacket,         --          .startofpacket
			sink4_endofpacket    => crosser_016_out_endofpacket,           --          .endofpacket
			sink5_ready          => crosser_018_out_ready,                 --     sink5.ready
			sink5_valid          => crosser_018_out_valid,                 --          .valid
			sink5_channel        => crosser_018_out_channel,               --          .channel
			sink5_data           => crosser_018_out_data,                  --          .data
			sink5_startofpacket  => crosser_018_out_startofpacket,         --          .startofpacket
			sink5_endofpacket    => crosser_018_out_endofpacket,           --          .endofpacket
			sink6_ready          => crosser_020_out_ready,                 --     sink6.ready
			sink6_valid          => crosser_020_out_valid,                 --          .valid
			sink6_channel        => crosser_020_out_channel,               --          .channel
			sink6_data           => crosser_020_out_data,                  --          .data
			sink6_startofpacket  => crosser_020_out_startofpacket,         --          .startofpacket
			sink6_endofpacket    => crosser_020_out_endofpacket,           --          .endofpacket
			sink7_ready          => crosser_022_out_ready,                 --     sink7.ready
			sink7_valid          => crosser_022_out_valid,                 --          .valid
			sink7_channel        => crosser_022_out_channel,               --          .channel
			sink7_data           => crosser_022_out_data,                  --          .data
			sink7_startofpacket  => crosser_022_out_startofpacket,         --          .startofpacket
			sink7_endofpacket    => crosser_022_out_endofpacket,           --          .endofpacket
			sink8_ready          => crosser_024_out_ready,                 --     sink8.ready
			sink8_valid          => crosser_024_out_valid,                 --          .valid
			sink8_channel        => crosser_024_out_channel,               --          .channel
			sink8_data           => crosser_024_out_data,                  --          .data
			sink8_startofpacket  => crosser_024_out_startofpacket,         --          .startofpacket
			sink8_endofpacket    => crosser_024_out_endofpacket,           --          .endofpacket
			sink9_ready          => width_adapter_003_src_ready,           --     sink9.ready
			sink9_valid          => width_adapter_003_src_valid,           --          .valid
			sink9_channel        => width_adapter_003_src_channel,         --          .channel
			sink9_data           => width_adapter_003_src_data,            --          .data
			sink9_startofpacket  => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink9_endofpacket    => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink10_ready         => crosser_026_out_ready,                 --    sink10.ready
			sink10_valid         => crosser_026_out_valid,                 --          .valid
			sink10_channel       => crosser_026_out_channel,               --          .channel
			sink10_data          => crosser_026_out_data,                  --          .data
			sink10_startofpacket => crosser_026_out_startofpacket,         --          .startofpacket
			sink10_endofpacket   => crosser_026_out_endofpacket,           --          .endofpacket
			sink11_ready         => crosser_028_out_ready,                 --    sink11.ready
			sink11_valid         => crosser_028_out_valid,                 --          .valid
			sink11_channel       => crosser_028_out_channel,               --          .channel
			sink11_data          => crosser_028_out_data,                  --          .data
			sink11_startofpacket => crosser_028_out_startofpacket,         --          .startofpacket
			sink11_endofpacket   => crosser_028_out_endofpacket            --          .endofpacket
		);

	rsp_xbar_mux_002 : component DE4_QSYS_rsp_xbar_mux_002
		port map (
			clk                 => mem_if_ddr2_emif_afi_clk_clk,       --       clk.clk
			reset               => rst_controller_reset_out_reset,     -- clk_reset.reset
			src_ready           => rsp_xbar_mux_002_src_ready,         --       src.ready
			src_valid           => rsp_xbar_mux_002_src_valid,         --          .valid
			src_data            => rsp_xbar_mux_002_src_data,          --          .data
			src_channel         => rsp_xbar_mux_002_src_channel,       --          .channel
			src_startofpacket   => rsp_xbar_mux_002_src_startofpacket, --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_002_src_endofpacket,   --          .endofpacket
			sink0_ready         => crosser_017_out_ready,              --     sink0.ready
			sink0_valid         => crosser_017_out_valid,              --          .valid
			sink0_channel       => crosser_017_out_channel,            --          .channel
			sink0_data          => crosser_017_out_data,               --          .data
			sink0_startofpacket => crosser_017_out_startofpacket,      --          .startofpacket
			sink0_endofpacket   => crosser_017_out_endofpacket,        --          .endofpacket
			sink1_ready         => crosser_019_out_ready,              --     sink1.ready
			sink1_valid         => crosser_019_out_valid,              --          .valid
			sink1_channel       => crosser_019_out_channel,            --          .channel
			sink1_data          => crosser_019_out_data,               --          .data
			sink1_startofpacket => crosser_019_out_startofpacket,      --          .startofpacket
			sink1_endofpacket   => crosser_019_out_endofpacket,        --          .endofpacket
			sink2_ready         => crosser_021_out_ready,              --     sink2.ready
			sink2_valid         => crosser_021_out_valid,              --          .valid
			sink2_channel       => crosser_021_out_channel,            --          .channel
			sink2_data          => crosser_021_out_data,               --          .data
			sink2_startofpacket => crosser_021_out_startofpacket,      --          .startofpacket
			sink2_endofpacket   => crosser_021_out_endofpacket,        --          .endofpacket
			sink3_ready         => crosser_023_out_ready,              --     sink3.ready
			sink3_valid         => crosser_023_out_valid,              --          .valid
			sink3_channel       => crosser_023_out_channel,            --          .channel
			sink3_data          => crosser_023_out_data,               --          .data
			sink3_startofpacket => crosser_023_out_startofpacket,      --          .startofpacket
			sink3_endofpacket   => crosser_023_out_endofpacket,        --          .endofpacket
			sink4_ready         => crosser_025_out_ready,              --     sink4.ready
			sink4_valid         => crosser_025_out_valid,              --          .valid
			sink4_channel       => crosser_025_out_channel,            --          .channel
			sink4_data          => crosser_025_out_data,               --          .data
			sink4_startofpacket => crosser_025_out_startofpacket,      --          .startofpacket
			sink4_endofpacket   => crosser_025_out_endofpacket,        --          .endofpacket
			sink5_ready         => crosser_027_out_ready,              --     sink5.ready
			sink5_valid         => crosser_027_out_valid,              --          .valid
			sink5_channel       => crosser_027_out_channel,            --          .channel
			sink5_data          => crosser_027_out_data,               --          .data
			sink5_startofpacket => crosser_027_out_startofpacket,      --          .startofpacket
			sink5_endofpacket   => crosser_027_out_endofpacket,        --          .endofpacket
			sink6_ready         => crosser_029_out_ready,              --     sink6.ready
			sink6_valid         => crosser_029_out_valid,              --          .valid
			sink6_channel       => crosser_029_out_channel,            --          .channel
			sink6_data          => crosser_029_out_data,               --          .data
			sink6_startofpacket => crosser_029_out_startofpacket,      --          .startofpacket
			sink6_endofpacket   => crosser_029_out_endofpacket         --          .endofpacket
		);

	width_adapter : component DE4_QSYS_width_adapter
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset             => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid          => cmd_xbar_demux_001_src9_valid,         --      sink.valid
			in_channel        => cmd_xbar_demux_001_src9_channel,       --          .channel
			in_startofpacket  => cmd_xbar_demux_001_src9_startofpacket, --          .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,   --          .endofpacket
			in_ready          => cmd_xbar_demux_001_src9_ready,         --          .ready
			in_data           => cmd_xbar_demux_001_src9_data,          --          .data
			out_endofpacket   => width_adapter_src_endofpacket,         --       src.endofpacket
			out_data          => width_adapter_src_data,                --          .data
			out_channel       => width_adapter_src_channel,             --          .channel
			out_valid         => width_adapter_src_valid,               --          .valid
			out_ready         => width_adapter_src_ready,               --          .ready
			out_startofpacket => width_adapter_src_startofpacket        --          .startofpacket
		);

	width_adapter_001 : component DE4_QSYS_width_adapter
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset             => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid          => cmd_xbar_demux_003_src0_valid,         --      sink.valid
			in_channel        => cmd_xbar_demux_003_src0_channel,       --          .channel
			in_startofpacket  => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			in_endofpacket    => cmd_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			in_ready          => cmd_xbar_demux_003_src0_ready,         --          .ready
			in_data           => cmd_xbar_demux_003_src0_data,          --          .data
			out_endofpacket   => width_adapter_001_src_endofpacket,     --       src.endofpacket
			out_data          => width_adapter_001_src_data,            --          .data
			out_channel       => width_adapter_001_src_channel,         --          .channel
			out_valid         => width_adapter_001_src_valid,           --          .valid
			out_ready         => width_adapter_001_src_ready,           --          .ready
			out_startofpacket => width_adapter_001_src_startofpacket    --          .startofpacket
		);

	width_adapter_002 : component DE4_QSYS_width_adapter_002
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset             => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid          => cmd_xbar_demux_004_src0_valid,         --      sink.valid
			in_channel        => cmd_xbar_demux_004_src0_channel,       --          .channel
			in_startofpacket  => cmd_xbar_demux_004_src0_startofpacket, --          .startofpacket
			in_endofpacket    => cmd_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			in_ready          => cmd_xbar_demux_004_src0_ready,         --          .ready
			in_data           => cmd_xbar_demux_004_src0_data,          --          .data
			out_endofpacket   => width_adapter_002_src_endofpacket,     --       src.endofpacket
			out_data          => width_adapter_002_src_data,            --          .data
			out_channel       => width_adapter_002_src_channel,         --          .channel
			out_valid         => width_adapter_002_src_valid,           --          .valid
			out_ready         => width_adapter_002_src_ready,           --          .ready
			out_startofpacket => width_adapter_002_src_startofpacket    --          .startofpacket
		);

	width_adapter_003 : component DE4_QSYS_width_adapter_003
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset             => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			in_valid          => rsp_xbar_demux_009_src0_valid,         --      sink.valid
			in_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			in_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			in_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			in_ready          => rsp_xbar_demux_009_src0_ready,         --          .ready
			in_data           => rsp_xbar_demux_009_src0_data,          --          .data
			out_endofpacket   => width_adapter_003_src_endofpacket,     --       src.endofpacket
			out_data          => width_adapter_003_src_data,            --          .data
			out_channel       => width_adapter_003_src_channel,         --          .channel
			out_valid         => width_adapter_003_src_valid,           --          .valid
			out_ready         => width_adapter_003_src_ready,           --          .ready
			out_startofpacket => width_adapter_003_src_startofpacket    --          .startofpacket
		);

	width_adapter_004 : component DE4_QSYS_width_adapter_003
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset             => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			in_valid          => rsp_xbar_demux_009_src1_valid,         --      sink.valid
			in_channel        => rsp_xbar_demux_009_src1_channel,       --          .channel
			in_startofpacket  => rsp_xbar_demux_009_src1_startofpacket, --          .startofpacket
			in_endofpacket    => rsp_xbar_demux_009_src1_endofpacket,   --          .endofpacket
			in_ready          => rsp_xbar_demux_009_src1_ready,         --          .ready
			in_data           => rsp_xbar_demux_009_src1_data,          --          .data
			out_endofpacket   => width_adapter_004_src_endofpacket,     --       src.endofpacket
			out_data          => width_adapter_004_src_data,            --          .data
			out_channel       => width_adapter_004_src_channel,         --          .channel
			out_valid         => width_adapter_004_src_valid,           --          .valid
			out_ready         => width_adapter_004_src_ready,           --          .ready
			out_startofpacket => width_adapter_004_src_startofpacket    --          .startofpacket
		);

	width_adapter_005 : component DE4_QSYS_width_adapter_005
		port map (
			clk               => mem_if_ddr2_emif_afi_clk_clk,          --       clk.clk
			reset             => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			in_valid          => rsp_xbar_demux_009_src2_valid,         --      sink.valid
			in_channel        => rsp_xbar_demux_009_src2_channel,       --          .channel
			in_startofpacket  => rsp_xbar_demux_009_src2_startofpacket, --          .startofpacket
			in_endofpacket    => rsp_xbar_demux_009_src2_endofpacket,   --          .endofpacket
			in_ready          => rsp_xbar_demux_009_src2_ready,         --          .ready
			in_data           => rsp_xbar_demux_009_src2_data,          --          .data
			out_endofpacket   => width_adapter_005_src_endofpacket,     --       src.endofpacket
			out_data          => width_adapter_005_src_data,            --          .data
			out_channel       => width_adapter_005_src_channel,         --          .channel
			out_valid         => width_adapter_005_src_valid,           --          .valid
			out_ready         => width_adapter_005_src_ready,           --          .ready
			out_startofpacket => width_adapter_005_src_startofpacket    --          .startofpacket
		);

	crosser : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src3_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src3_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src3_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src3_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src3_data,          --              .data
			out_ready         => crosser_out_ready,                     --           out.ready
			out_valid         => crosser_out_valid,                     --              .valid
			out_startofpacket => crosser_out_startofpacket,             --              .startofpacket
			out_endofpacket   => crosser_out_endofpacket,               --              .endofpacket
			out_channel       => crosser_out_channel,                   --              .channel
			out_data          => crosser_out_data                       --              .data
		);

	crosser_001 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src4_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src4_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src4_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src4_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src4_data,          --              .data
			out_ready         => crosser_001_out_ready,                 --           out.ready
			out_valid         => crosser_001_out_valid,                 --              .valid
			out_startofpacket => crosser_001_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_001_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_001_out_channel,               --              .channel
			out_data          => crosser_001_out_data                   --              .data
		);

	crosser_002 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src5_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src5_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src5_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src5_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src5_data,          --              .data
			out_ready         => crosser_002_out_ready,                 --           out.ready
			out_valid         => crosser_002_out_valid,                 --              .valid
			out_startofpacket => crosser_002_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_002_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_002_out_channel,               --              .channel
			out_data          => crosser_002_out_data                   --              .data
		);

	crosser_003 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src6_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src6_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src6_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src6_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src6_data,          --              .data
			out_ready         => crosser_003_out_ready,                 --           out.ready
			out_valid         => crosser_003_out_valid,                 --              .valid
			out_startofpacket => crosser_003_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_003_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_003_out_channel,               --              .channel
			out_data          => crosser_003_out_data                   --              .data
		);

	crosser_004 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src7_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src7_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src7_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src7_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src7_data,          --              .data
			out_ready         => crosser_004_out_ready,                 --           out.ready
			out_valid         => crosser_004_out_valid,                 --              .valid
			out_startofpacket => crosser_004_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_004_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_004_out_channel,               --              .channel
			out_data          => crosser_004_out_data                   --              .data
		);

	crosser_005 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src8_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src8_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src8_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src8_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src8_data,          --              .data
			out_ready         => crosser_005_out_ready,                 --           out.ready
			out_valid         => crosser_005_out_valid,                 --              .valid
			out_startofpacket => crosser_005_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_005_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_005_out_channel,               --              .channel
			out_data          => crosser_005_out_data                   --              .data
		);

	crosser_006 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,           --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,         --  in_clk_reset.reset
			out_clk           => clk_clk,                                --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,     -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src10_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src10_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src10_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src10_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src10_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src10_data,          --              .data
			out_ready         => crosser_006_out_ready,                  --           out.ready
			out_valid         => crosser_006_out_valid,                  --              .valid
			out_startofpacket => crosser_006_out_startofpacket,          --              .startofpacket
			out_endofpacket   => crosser_006_out_endofpacket,            --              .endofpacket
			out_channel       => crosser_006_out_channel,                --              .channel
			out_data          => crosser_006_out_data                    --              .data
		);

	crosser_007 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,           --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,         --  in_clk_reset.reset
			out_clk           => clk_clk,                                --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,     -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src11_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src11_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src11_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src11_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src11_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src11_data,          --              .data
			out_ready         => crosser_007_out_ready,                  --           out.ready
			out_valid         => crosser_007_out_valid,                  --              .valid
			out_startofpacket => crosser_007_out_startofpacket,          --              .startofpacket
			out_endofpacket   => crosser_007_out_endofpacket,            --              .endofpacket
			out_channel       => crosser_007_out_channel,                --              .channel
			out_data          => crosser_007_out_data                    --              .data
		);

	crosser_008 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src0_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src0_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src0_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src0_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src0_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src0_data,          --              .data
			out_ready         => crosser_008_out_ready,                 --           out.ready
			out_valid         => crosser_008_out_valid,                 --              .valid
			out_startofpacket => crosser_008_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_008_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_008_out_channel,               --              .channel
			out_data          => crosser_008_out_data                   --              .data
		);

	crosser_009 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src1_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src1_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src1_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src1_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src1_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src1_data,          --              .data
			out_ready         => crosser_009_out_ready,                 --           out.ready
			out_valid         => crosser_009_out_valid,                 --              .valid
			out_startofpacket => crosser_009_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_009_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_009_out_channel,               --              .channel
			out_data          => crosser_009_out_data                   --              .data
		);

	crosser_010 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src2_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src2_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src2_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src2_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src2_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src2_data,          --              .data
			out_ready         => crosser_010_out_ready,                 --           out.ready
			out_valid         => crosser_010_out_valid,                 --              .valid
			out_startofpacket => crosser_010_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_010_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_010_out_channel,               --              .channel
			out_data          => crosser_010_out_data                   --              .data
		);

	crosser_011 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src3_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src3_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src3_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src3_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src3_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src3_data,          --              .data
			out_ready         => crosser_011_out_ready,                 --           out.ready
			out_valid         => crosser_011_out_valid,                 --              .valid
			out_startofpacket => crosser_011_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_011_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_011_out_channel,               --              .channel
			out_data          => crosser_011_out_data                   --              .data
		);

	crosser_012 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src4_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src4_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src4_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src4_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src4_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src4_data,          --              .data
			out_ready         => crosser_012_out_ready,                 --           out.ready
			out_valid         => crosser_012_out_valid,                 --              .valid
			out_startofpacket => crosser_012_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_012_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_012_out_channel,               --              .channel
			out_data          => crosser_012_out_data                   --              .data
		);

	crosser_013 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src5_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src5_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src5_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src5_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src5_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src5_data,          --              .data
			out_ready         => crosser_013_out_ready,                 --           out.ready
			out_valid         => crosser_013_out_valid,                 --              .valid
			out_startofpacket => crosser_013_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_013_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_013_out_channel,               --              .channel
			out_data          => crosser_013_out_data                   --              .data
		);

	crosser_014 : component DE4_QSYS_crosser
		port map (
			in_clk            => mem_if_ddr2_emif_afi_clk_clk,          --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src6_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src6_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src6_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src6_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src6_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src6_data,          --              .data
			out_ready         => crosser_014_out_ready,                 --           out.ready
			out_valid         => crosser_014_out_valid,                 --              .valid
			out_startofpacket => crosser_014_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_014_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_014_out_channel,               --              .channel
			out_data          => crosser_014_out_data                   --              .data
		);

	crosser_015 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_003_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_003_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_003_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_003_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_003_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_003_src0_data,          --              .data
			out_ready         => crosser_015_out_ready,                 --           out.ready
			out_valid         => crosser_015_out_valid,                 --              .valid
			out_startofpacket => crosser_015_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_015_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_015_out_channel,               --              .channel
			out_data          => crosser_015_out_data                   --              .data
		);

	crosser_016 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_004_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_004_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_004_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_004_src0_data,          --              .data
			out_ready         => crosser_016_out_ready,                 --           out.ready
			out_valid         => crosser_016_out_valid,                 --              .valid
			out_startofpacket => crosser_016_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_016_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_016_out_channel,               --              .channel
			out_data          => crosser_016_out_data                   --              .data
		);

	crosser_017 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_004_src1_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_004_src1_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_004_src1_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_004_src1_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_004_src1_channel,       --              .channel
			in_data           => rsp_xbar_demux_004_src1_data,          --              .data
			out_ready         => crosser_017_out_ready,                 --           out.ready
			out_valid         => crosser_017_out_valid,                 --              .valid
			out_startofpacket => crosser_017_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_017_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_017_out_channel,               --              .channel
			out_data          => crosser_017_out_data                   --              .data
		);

	crosser_018 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_005_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_005_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_005_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_005_src0_data,          --              .data
			out_ready         => crosser_018_out_ready,                 --           out.ready
			out_valid         => crosser_018_out_valid,                 --              .valid
			out_startofpacket => crosser_018_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_018_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_018_out_channel,               --              .channel
			out_data          => crosser_018_out_data                   --              .data
		);

	crosser_019 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_005_src1_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_005_src1_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_005_src1_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_005_src1_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_005_src1_channel,       --              .channel
			in_data           => rsp_xbar_demux_005_src1_data,          --              .data
			out_ready         => crosser_019_out_ready,                 --           out.ready
			out_valid         => crosser_019_out_valid,                 --              .valid
			out_startofpacket => crosser_019_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_019_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_019_out_channel,               --              .channel
			out_data          => crosser_019_out_data                   --              .data
		);

	crosser_020 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_006_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_006_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_006_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_006_src0_data,          --              .data
			out_ready         => crosser_020_out_ready,                 --           out.ready
			out_valid         => crosser_020_out_valid,                 --              .valid
			out_startofpacket => crosser_020_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_020_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_020_out_channel,               --              .channel
			out_data          => crosser_020_out_data                   --              .data
		);

	crosser_021 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_006_src1_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_006_src1_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_006_src1_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_006_src1_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_006_src1_channel,       --              .channel
			in_data           => rsp_xbar_demux_006_src1_data,          --              .data
			out_ready         => crosser_021_out_ready,                 --           out.ready
			out_valid         => crosser_021_out_valid,                 --              .valid
			out_startofpacket => crosser_021_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_021_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_021_out_channel,               --              .channel
			out_data          => crosser_021_out_data                   --              .data
		);

	crosser_022 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_007_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_007_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_007_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_007_src0_data,          --              .data
			out_ready         => crosser_022_out_ready,                 --           out.ready
			out_valid         => crosser_022_out_valid,                 --              .valid
			out_startofpacket => crosser_022_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_022_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_022_out_channel,               --              .channel
			out_data          => crosser_022_out_data                   --              .data
		);

	crosser_023 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_007_src1_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_007_src1_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_007_src1_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_007_src1_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_007_src1_channel,       --              .channel
			in_data           => rsp_xbar_demux_007_src1_data,          --              .data
			out_ready         => crosser_023_out_ready,                 --           out.ready
			out_valid         => crosser_023_out_valid,                 --              .valid
			out_startofpacket => crosser_023_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_023_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_023_out_channel,               --              .channel
			out_data          => crosser_023_out_data                   --              .data
		);

	crosser_024 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_008_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_008_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_008_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_008_src0_data,          --              .data
			out_ready         => crosser_024_out_ready,                 --           out.ready
			out_valid         => crosser_024_out_valid,                 --              .valid
			out_startofpacket => crosser_024_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_024_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_024_out_channel,               --              .channel
			out_data          => crosser_024_out_data                   --              .data
		);

	crosser_025 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_008_src1_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_008_src1_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_008_src1_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_008_src1_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_008_src1_channel,       --              .channel
			in_data           => rsp_xbar_demux_008_src1_data,          --              .data
			out_ready         => crosser_025_out_ready,                 --           out.ready
			out_valid         => crosser_025_out_valid,                 --              .valid
			out_startofpacket => crosser_025_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_025_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_025_out_channel,               --              .channel
			out_data          => crosser_025_out_data                   --              .data
		);

	crosser_026 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_010_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_010_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_010_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_010_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_010_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_010_src0_data,          --              .data
			out_ready         => crosser_026_out_ready,                 --           out.ready
			out_valid         => crosser_026_out_valid,                 --              .valid
			out_startofpacket => crosser_026_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_026_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_026_out_channel,               --              .channel
			out_data          => crosser_026_out_data                   --              .data
		);

	crosser_027 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_010_src1_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_010_src1_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_010_src1_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_010_src1_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_010_src1_channel,       --              .channel
			in_data           => rsp_xbar_demux_010_src1_data,          --              .data
			out_ready         => crosser_027_out_ready,                 --           out.ready
			out_valid         => crosser_027_out_valid,                 --              .valid
			out_startofpacket => crosser_027_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_027_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_027_out_channel,               --              .channel
			out_data          => crosser_027_out_data                   --              .data
		);

	crosser_028 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_011_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_011_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_011_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_011_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_011_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_011_src0_data,          --              .data
			out_ready         => crosser_028_out_ready,                 --           out.ready
			out_valid         => crosser_028_out_valid,                 --              .valid
			out_startofpacket => crosser_028_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_028_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_028_out_channel,               --              .channel
			out_data          => crosser_028_out_data                   --              .data
		);

	crosser_029 : component DE4_QSYS_crosser
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => mem_if_ddr2_emif_afi_clk_clk,          --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_011_src1_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_011_src1_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_011_src1_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_011_src1_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_011_src1_channel,       --              .channel
			in_data           => rsp_xbar_demux_011_src1_data,          --              .data
			out_ready         => crosser_029_out_ready,                 --           out.ready
			out_valid         => crosser_029_out_valid,                 --              .valid
			out_startofpacket => crosser_029_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_029_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_029_out_channel,               --              .channel
			out_data          => crosser_029_out_data                   --              .data
		);

	irq_mapper : component DE4_QSYS_irq_mapper
		port map (
			clk           => mem_if_ddr2_emif_afi_clk_clk,   --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_qsys_d_irq_irq            --    sender.irq
		);

	irq_synchronizer : component DE4_QSYS_irq_synchronizer
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => mem_if_ddr2_emif_afi_clk_clk,       --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	irq_synchronizer_001 : component DE4_QSYS_irq_synchronizer
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => mem_if_ddr2_emif_afi_clk_clk,       --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	irq_synchronizer_002 : component DE4_QSYS_irq_synchronizer
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => mem_if_ddr2_emif_afi_clk_clk,       --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver3_irq            --             sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	led_s1_translator_avalon_anti_slave_0_write_ports_inv <= not led_s1_translator_avalon_anti_slave_0_write;

	timer_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_s1_translator_avalon_anti_slave_0_write;

	spi_2_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv <= not spi_2_spi_control_port_translator_avalon_anti_slave_0_write;

	spi_2_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv <= not spi_2_spi_control_port_translator_avalon_anti_slave_0_read;

	mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_inv <= not mem_if_ddr2_emif_avl_waitrequest;

	spi_1_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv <= not spi_1_spi_control_port_translator_avalon_anti_slave_0_write;

	spi_1_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv <= not spi_1_spi_control_port_translator_avalon_anti_slave_0_read;

	no_of_cam_channels_s1_translator_avalon_anti_slave_0_write_ports_inv <= not no_of_cam_channels_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	mem_if_ddr2_emif_afi_reset_reset_ports_inv <= not mem_if_ddr2_emif_afi_reset_reset;

end architecture rtl; -- of DE4_QSYS
