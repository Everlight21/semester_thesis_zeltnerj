��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X������]u�.���\�KI�?�5Z�>�%i�v!����wkhO�������X{�ٸ��Tb� )C(���B��r��q��T}��4�I�����#U�����Q�[Z'��~�����T�D��[�U8g���T�(��QƘ︟��^�������3e��,���	�q�W��e�P�����y���	����'s'��%n7	�/%Ӫ�{�����cpW]�+�E��SC��v�ɂ�)ٗ�u�#Z�ޢ?;C���ɚ�=�2f"{vZ����-q&� �Vr`�hs��e�<��#���>�OMx�g���A?'���M���Ҥ���7Zι.�ݷ�:���vZa�9��)$����&��^�-; ��B=g�<2�Zu�S��4���~�20~���Oi�����;���()�%6�J����n�C���z������O[Q�j�%����e��r1��#Uu�g^(��(��x\I�;�m�(��"[�m��r� �xk<�4��8l�1f�Q!�B���5+fa��&
x�R�J���Ku�o��(�gp��C籿砢X����}�`����\�=o����;ǘҨK�L9�!!AS�Ϯ�I\\Q�ΈYI����	�Y��@
��Q���+�0��ǁ��^�o��z�bV�k&�\�hLX�
��R��#�����c_ma�[��
0���9�O�����)��c2u��Q�����b�]�'-�����|�M/� �t�h��=UU�o�='I�$|
���ܷ�\�w�jD���Z���*��^_�>W%��@RK9EFg,i���,A��=f:UͲ�v1֟�.&�]QÝ��j�(&8�7���*�6�t4�K;��9�u��a25s�$��^�r�P����I����g�U؀�T1��b�y���#OW�9��Wע�����b�����2�c-7E���������hv�,t�$1�"!��nu�����<�=Ͼ�����8��w[q�ϛ(�_%���P8�ԍe��	澢O���J\�.�����.�K{��t�~�'$�{�<ho�gC������	[�N����01�ɘ�1K�Slk�'͎a��t�$���i����w8�ml��m������n��!�g���k�+�=��Q��mt�CSVȮ��S�;�,�aH9�� /wֽ�\(��qw�(F�B��I>��9z��n��~>��jiĿ�-��+��4qКfoE���n[_&�v�)����xL�M	�x|��-�Zv�&Գ���^�ƞX=���S���/��J:����J��o*0���f{J�X�0�B��Nn6
翊���=|�>W�����C,g,P�lw�jq��0�̏A��2������6�D�x`0>�^�{n������Z�_��h��9�fINa�a���.	�:6t�'��+Â3�"B��q ΧW����	L�����"D������ė$�I!~I"����� �SS�݁� ����g�~j�̍��X#�;�\���#+�!6�&R��e�7��.9��4����۷5uk��e֕�J�Ba����_�<�k׆τ1�����d�K���|L��%Sv_o�_^�=�K�2
��ϖ.��֨���wI(:�&��kg_�e��r\	�
A����&gox��VnA�sI2�<X0�	�WH�[�X?"k�G�$&jb[�������M9����Օ:�GX���/]Q|txo~i�9� B� ���9hW����`L��q�a��v_�7<��r$E�n�vl���2y>�]�4��L�a�����|n���#1��:��S}d���ӿA
W�.޲+��L���+ʏY(%�D�爏�^�S��2v�H0��JC���|��y\7�1xR$-�5/���8�!3�&�c�z����_�<��~��b��Y��lG2�E}S�,QjƼJ�n��vy�bt�P�������-[��θ5�+�p�����y���C�ReY��O�L2�N�m��Y��/�����g��u�6�z�����u�P7p5ϫ��Z�3��v�{����\��4�-�bs9lI5y�xBo�mC�]�<M#jלn��5ElU���p�,�}l�e$z������o�����9~�]�!�%��I�� [�Q�	��J^0@�K����\T����8úHB3��ej�b #��o�����~A�A���XZV�O�����$v�&���/Yd{՚��*H���K�o$��F�iMi�Hȓ3^z7�6��;w_����4oCػ�tP ���0h7{��KP��ge�����f1�Yy/�XѫM.z���X��#��{ܲZHz�H\m%���R�g��岖:�i�L�8n	QN�>�z�p���;u����W�TrmPS�c�l&ןt��y��rp�j6z�ry#�T�N���n��j�[|!�-��}�3h���;L���!ry��p�0ϩ��"^��DA�j����i��\�+X �)`�6BNÃ�B�ag`ct�q��ƴ,͉�s�
>�� (���U�Yt;���`$�>2�	�������W���v�T��ݿ�p��t���;	_
�t�);� rӞ�ɸ˖@�(����<�'���,�����ڭW��HD����q+���Z�㮫=g�� N_v8�Am>�%;��9F�W��[O�a���W��ꆻj���˶�W
-��u�(�1ۀp+hH���c�
6�wՀ�m���"n�!��s=��v��*w|��$͗�ʢ��O>�;��]Q+J.��SC�U��I%�n>��Q�@��ǭZB��Y�^�G��p�ݬ�b���9G��<hs��n	�kQ��Nq��y�~s)�26d43c�y��R[�)�'gL
����	��\?���VY�}~_��*'$�S��5���z_�H]�H5
o��gV�{��b5�dY{�I�z��z�E�1��� �l�=��1��в��s����%`b�3<�VD���o�?�挂Ae�w���&f�/	�E.���_ޝ����*�E���/��][����i@G�)�li����%!��z�=��񁣛�*�Sz?iNk/�Q�W�b�e�E��Q�H�^�ϗ4���>D�����*�����v´Ӵ�u私�Q���g9��kHL���Ā�n}(�	<��8�2��5M��d�U:$�|T&�>�"7i�����G����FI��3�4�*��6�Q����&-�U-K�<�a�|�$��ˎB��B8�N��s�&���P�1�k�e�̦��aQ��I�GT,�7[��r��S�M�/�����.��Z��y�H�/OK�'f���O��B`%3���i7y"ӵ%�%�}����kZn��DM�t ���BJDl���"CA�a
87��et�9{�P�+�6������r�(��ۺ�L��Ŕ���k#>:~�^	�3���T��<-��E	��+M���Uj�i׮�KlU�'�AU�~:��3���uU��Ō�����n���\S���ʩ	~µ�А-��1����(
+Ԝ!^����3Z��+�D-���?��ލ�1�Z%S���7�	�̮Sl���O��U���N�L	koUq����T��Q.�s��������q�`E�rW��	�"G<ٚۉ̬G9{9����Y���@�������	��9�U����� �ˉ�I��[CM�Щ;K�7`˖M���Ƃ������8�!J$Vٲ��#���u�)��FX=�����_z��F*YZ�x�y9�#ٔߚQ�fj��'"�sD�]��:�څs���ۭ�~�X���'��Ϝ%d�u���gu$)R���i~��9[��n�������2uo?R*T�x5�g7#��U�U� ҁg�*�\�F�BB�HU�x1rJgŲ���=�gjl�V6��
e�f��ʯ�+D���g9	���[��<5��v�F,)� NV��<\��$�S���jU�!eO�_�0ې�b������!Jk�at��|�j����u�B[�ڎ�M�zW_���O���YOKh6*
H`@}M��@�����'@g���!fa�]�K����u� j������ۡ��rB)�C�ٮ:��u"R��	�a�=W���dY�
W� ���3w�Q�W��r'�Z}�[��b���%�v���!�\�Hn=��QzH.��D����v�YR"��a��Tv��S?��*���}�sr	��7f�S���f�/�
j��/�^�ڇ�.��&(�w��]��B5���-J�0��@���S�L�u�f(��z���Ïѡ���# �1���Aa��Ġ�AU* W���m ,z�T����}�\�I��o����n��6�2��^M�ц����}+����z#����������`��� G4�9�;0�T]ٷ � tj[IL���Ay�'x.��� ��V��`���McA�۝A��~��h�A��^�:�����:�>Ƅ8}��jY����Pb�Z�r��)�D��=�T��t�auRJ;t�b#x��KZ���_"����$Z��e��ԟ@�d\�obƢ�݂pb�gk����.͐��[�dl�А��݅��Z�������f_d�ή9z�m"�M @�Șp�+d�z�hצ�� _�1#�(��+�OP3wCj,������pEv�1���iPT�9�;�L�ůEId7�dz��Ui�bL^��6��fu)U\����%i�z��l������t�ě �� 0B�7�k?t�qK}R���,�q���3��d�����n�ýz�-�Po���Zw} �<��D��x0B�v4�Ĉ�%���T4��Ƀ�fe�/M1a�[����$Ԇ-�9�//Vj�K�q��������WGڢ`:��/�-���
Ųd��G���f�M��S�9P���T�%���3`�䕭�-�JD��7գm]�����cF�n�g���56#�e���4mB\����g�${�zV���D���9��������ҩ�\�g��ЊAC��"�h	�Do2z�"��kQ��9W|�*�k�J��H���ǩ�Ȭ��Hb}H{����Y�f��=�=�=�\ч(2��B��>ɮ��ٟ�5Y��-!ɉ#���_�I����WMK��4U	����@<�n�
b.��H-s�ķ:Qe?�+���6̦�Y�p�ێ���]!�� |(3��{����~���V�#غ�dM������.�ϊ�;���o����Y��G��*H��3��1�=9\���=�s{�ln�lt�P����+~؞��u�7=�y1��^��1�3�ꙛQ� ��%n��v/y�Id(yXA�E� ��O���S��2F�/Z"����F�\�����m?Y|��p?�PG��=j��fqF$I��E��nX�v�]��!~���YF].��b5�nq��;��D�s�p]�l*\V�lS�-�����5;=��,� x͂�a�����%,�w(w��[���6��磻p��{��ǔ���I�KIC�t?e+��m�ʩ���K&�	�{����w򖢻���]h 	�lՒd�)9����r�)| ,���h3�Y��_�-~%�s��U\���AZI.?H�We�?K��:6�[�,��T��"s�~:�� ����.G���"�7�a��	�J9�5(��)�a���\���}
Ժ����5%�ڋN�ey��;��Õ�v"��E��|�S����7ξ�&Ui*^�����\![�^"��]�)Gn
�f�r�B卶�j����$*��4wpQ-p��X����c������	RM/��$Rm%��0|�U�P��F�H/ܴ��kF߉.�G�#E�@j�02��ȉ�&1)!����� }��
���ke�7<N�e�-Z�޴�(�&6�[��3�ĊռԿh@�!a��Y��_�/iF�/��u�V��4�#	�zfvc4�A+�%��.`���t�#@�~�>P�����5�
C�MVnu<"�x��ve�V�� �A�ڊ[��v�3"	8A�}~4j��.S�I1�F��j�N`)���aw�O�+�]M��(a-�	TJ�Ie�=N�	&S� z�_Ɉ�?iU�T���b��c͈p��]c�d�� w�f�ˈ��;�:Dξg�=��~��QEW;<�OO���h 3���V���J�څX<?}%���`� ����c(p����|���ὄag�;�J<�/�g��̫�}�c��[�I���5���7e�bb|�U�ŷבZq��k̯�`|� �ԉ��K�����wD��t�j%�yL}n��&\~�����O�ܭ�����5�7�[ޤP�Ye���ks�f~��Y�:�vKP�8�����W���;���#R��r�|5�zw֞7�#t��B�Ěb7W�a:���ȇ�t"��뒠��mH��?Y�X�n���N$W39�Cf�]�"kt{E���$i`q6�]��6�j��ܖ����!��_
\��y�Ts����t;�qqf�,��q�s;���Z��As�;� �Ư�}�5�g����3��� �Q���G��fNG���TBwen!��U%R)���R���u���!��v��vEYi
�?�HP]��qI�)af��>Y���]��+tE���c|��,���i�<�5��m%�G����\TU�Pޯ��<ѻ������v^N�b��ٗD!3V$PΠD�׈�����>���vollm�� L 2��xa�]��C�&k�?���,=^]�݄o$�S�w����㠟�Īj�a� ⍧�����pHٓ����=���	�@�r&��uJ7�����h�QM2�YJ���;
ћ,�cK#]�&g�+: �R߁�m�>ppޮ�P߶��"�����Ef�lxY�c�>���Y�ԗ�}�������״���� V�G�]���Vu�k�ʸ�ݗ.��T�@NIߎP�[g��%��+z/�$���07�GH����蒱Qĸ�@^��g]r��(ᩞs���Y�!��Y�>O�9���T7;�c�����8��y�hn��ۓh�;��#�s������C�*y:W�C�_{bP='�~��N�H���;�" �Z�o*dE�v�B~:���,�{�r8��`�I9���v����u��F{`��m���qY����^�ѝ!f�FR�8ތt� �+���4zϊ$⃉�@,���>l��:l�	�-��0VF�U���'�Q���C�>V�-� �^��f߿W4�N)`:[��0�i�?S�n�*,��;]"����/��;h1,{��$�oC�R�sx�nMb�ᦨ3��o	��(a%%bO� �Fv>�O��Vs�J}�$�����1�7��e`C�L��e�k	���'EE�ǽ�f��������A2���3��N�y<�t��)��B�9��g�X��d�Ӱ>����� a7`�ߠ���.�	������rq��I�F�sK������fn,�z�V2���`�cYe�9U�.����j�Ҕ��$8���(��a�x���;i���"�HB]��ݭ��8�V�KE'�/����R0�Տyf���M9�C�D�`p����|� �F���^���yH������N\Ro������Ɋ��%(@�?wY�l`	��aWT�H�rD!pu%������%�3��.SJ
��uH.B�,���a��Š[{㮸�6Rkn-��h*ٲ� 3؍�u�ê�*��'Ub��f����4���C���t���2շ�����9%ܫ��U�|#V*�2%A���.��L09]���HQi)�<���O8g�զRM���6�Fz�-���swNa�<�"k׬)'8�O1�������:\��M�9c��l�e
q��ց���P�u	T �X�c�e0_�}�{�%|q�L�:z���z�V���ꂟT�;6�8}o)�����8��4z�:��7l�_h&\�1�����6Y�ՃN#���A=�.1�J ��a��)op&�wxsˏ?�zn�b}�Ww*̔2����=�$ST*.yzHD�a���cx���ݍ�q���Y�=���ؿ���1ٯ�v�-Yh����ѨL��'�Y��s�-Y���Jۉ���R5^�)�CAԳ*����0�e����2}�ƥ_�p.����́���|��=N��!!�� OQ��K���XW�$��)����uc��P��j�:nP�`�`4(�~h|?04"(92�l~�#�V�;xu����H 9���/�,7i_3���c�VY3�H���e����:3���Bz <o��=�eǭ͵�[��?R�B��'��<�f��{Z1Ĵ;O	;��3����VOm3ؙ	�<,�yd�z��֖����lAu�qå~��og ߥ:Nudʉ�
��Y��� �;�1��\�������zjiK���k�!��$��i�k�`��`�$�U�������'������o��$�R��,ɿ��H��w�G�h�f�<�g��QWr%G ��g�V˚D��Q�%o���-���H���<�?����5�����h'd��U�t����%fv��f��M��',�*(�^�a���	j�._N�A,NQ)Z��ֿ ,���Në���T�ý4�C�kf���av�����j�y;�,�d���'N��t�j�[�;u_9��i�_��ñ1�K���`��h�/�����@�?.�����k&K���h��Dm$��d�}'R<��0��oKe�$R`�\��NmFӋ�~�������l�"w������Ů�v9�A��yo%�NŹ���K��֍�Ji��K]��D��Vxx�)&�&��h��H�f�zj�m��E'��!��:�>*���-�15c?u��grT�QE�lz��L��CRO(��pZ�5�˱�.��`h`�@9jm���@ߠZ�� �Ȩ�td��R\�*��������Q����^�8S�om�ི���^N�j{���N
&�=]����O�8
 ׁ��]>��ćQ��&w�k�G��?Z���AUG_�:a�<��Ө�� o�V��Ôh������T�����Uǉ3N�m$n��ф5��d��\����!G���)�������&��'�����S
���X�<-��51����߭�ӑ[e��eU� �/ a���T��������Lؿ6J����?��5T �I$��;�jSW�	��7�r����͹�Q6�$����ٖ���������e>^����c�u%y��֗�t?#>H�R&��ΝIE�Z�Zmһ���b���n�i.>�B�7מu�C:�\X����x#"�T�4m��sIA���'��_փA U�׌��Ű"0�=,4���b��L�_�Է��m�rHN��S�*ꋻca�U뮿��t�0��;�����'':�K�!��B( ��	gd���2,�3Π$7�nJ���ν� \����ҙ4Q0:]�QϹEZ���������ln�Q�$��>�g�Z֌f��y���|��(���'e�.���Yխ��y��	R��m��K�z��y��B�����B�Z$J�Q=�Y��LW�O2��(tՉ�V��I-�g�_jH��!���A7�=s
ǌ���t��j"���L.!�:��F!�o��G�}H���,ߛ?[mK_������ர?S]I:k��cs!�x>��{4)���)��m�!G�/M��6�څI�)jX�I�B��,_��OV0cSY-�&𫼘kS��2(�Ph�̃ �jU-�.ڗ��B�bp+�� ���o��m�U�6
��|z��Uf��� �|V�c�U�����M��9�D�e�ނ��� ��'�%��"a��5��ݖ�׋2jͨw���}LI�=d"NT�W�Bix����97�¯�3<!���*nrs{������v�#&�}i+�`j�k-�:q��{O����l6~�!�ڗo8�F8��w!g.>\�6���u�� :��^0�n1<��VD�2��6��Rf��]�n�4At��D��w���
g�"�5��$��d:8;[1���.Y�A�B��?�g���U Ǉ�kN�v��\��*�Q���?�j3� ���Br��`���7��j�h�BB���)">��_��������0`í�Qe�KM�4(7���+��d�0��'<�a�2Z�K_���g�SX���i��A����.*�#���X`�;�X���D튼��U-D��)* ���aam�Of��3���Kߓ}q�c����4l�QW�qL'^����muE��UQ���d2���$ׁۓ�X�{r�G�O"��,5]ۍ�a���F���Gru����,~O�K��0�b���F&wF8�;`��M�ZR���>]���(���I����!?����c+�VL^z0Wٓ�]���]+�sٲ��ҳ>�jD!��[����3�ft_�ic��\����ެ�0���`0u�d|(e��.�P2S@��f5D��K�A]@�V!�-F����>���|֌�`�Fk��}��s�#�1�[�g*�����N�-���1_Ƽ�����@�#U��֦Ÿ�@� �����-�����W��=�`�)u/Ig�#�����F��2{���㤊;D��$�0���X�У��&_R|��y���n8n��zV�0�O9G��u;j}�g�r]V��� >S�𷞗�q�]��_�af,�����V�|O6���,����W��ERM|�K=���~��Ֆ���@�ɽD�~��}:{��ȞD����t'&�Yb�g���ߚ�)"?Ap���'�W���U\8$����:�r4�"�VJ�!A� ��K��b;�{͝I�3��v�F�E��+�7�$	�zǯ��C4��#�j4�e�&qwg�N�c�rsC˕[�G��{�%`�`ˠi�÷�@�����w7���OJ��!�G���1�ҷ��o`�w��j٩w�|�6�
��Y�Ȳ��AV&>ن�1�C�B�}/~T�P�y	R�ʲ��'�[w��Ǫ$��G����6'#u�3
Y��^�o��"6�.B���w$���V(�P����
/�K���S��EI��+p�4�G�bY�&%���K]���NOup�Ϲ�X�s���1�����R��ܻ�l'#ᏡR�i����~�jC*���e���g\�j�_>�:Ɋ�U�rÚ� 2&a���Q�z8zV��d�zw�8m6�.��4ۀ�@ؓ��?饞��@�o�T
.A$���Ӫ���z�޳'o�ᮣ�B�1�M�;'}�9xՄA��<j���^��f�ㆾ{����I أ7��F?Vu�Pt�u�%iu�5"��\�ߵ͆�6���ع�u[y7�7�F��'g�V4P�C�v�1`y�(|��W�{��~V�����B!I�DDf1oE��(�|�D�የ��	����4h �R�w#Qt��*�$za����@D�l@`����5F7]>���۫��ok�I�tU�j�i�����y[�s+��O�ti����)
 g4S;�[.+J�\ԫ��dWs�;��;^Ph�;�}o���O��!G�t�O�������dO����z����y��E?)� +l�{���Z�1I]汒�+��Cu=3E��jc.�oԽ�'��#�r�!�nnYą%���)V�����d���Qo аi��V���W��n�#-(xT	h�h=�~��v@>��~��-Sr�ʦ�E�=fgB�z�'�zX� `��x�ď�̺�mN}7��;p��e#�%��a��Y�+9��У/��g���`�4�T}{��-nQZ��p��KS$q���r�BG�
ZeMMQ��1��S1��؍�mt��T�%�I��pm�ê1�+t�'_����4�0M�Z��Zry3Y��7���\x�<�0��t���b#�{���ŤVk�N�qf}����5Ft�תyA��
��`��Ӆyc�xǵ�#4��,��_h�,��ɀ��7�\�n|�Xw�7����k��d��S׌�����&F���Jr��%�1�i�T�2��m�=��~R��5��'w�8��sӑuG�����u���f$�zlpx��ZHp}����p���J������
],�?ǲ"�V��+b�ipY?ip��Q �&���h�ҨOY�pq�&�v��W%jj�;/3�"ߥ5�ۮ]��d�?��pZ�M�ReH�᥾�#lCJ�A�,�N\�k�"gx��r��a�B��T{a�����=f�30d���
�,�8�x����?��U�\F�Όڪ���Iu��1Q\j�@u����Ө|�������ŴtMd_��k�a� 69��h/�U"B 8��{d�:��`y�t���(�����+5��G\X2�5��������R��s���i*Z��-1�*��٩O�\L�K�E��|�%r�,�a�^���	w���[�@�xUf!�>q>A���2ݜs��ue��Q@Uf��<�K�h�+M�X=�C8���#�������S�������Ov��r�$�xz����wQ��VE#.��b��TK�H���O�q�;�D��}$qr�i)^�hN��b���p���]}U�^�>����35ٝ�Xw���{th��wȴ���O=6#m!3m6��a�_)�����l��/�=�"-�N���#Lu��O�m�:zB;?6d���B>E?�����U%j�8l|mԼ>)�|G$ ����L3#����b��=�� s�	��5����c�b�l�9���]�(tD$���4�RI%@�}�g�e`�����T�x���Dϲ���������� r\�K;v�����X)�%�1\�K�)�O(��hU�+�4#�F��1�@ ȗ�!x�`2���/;�H;s�)���t��F{;��#6ү�����wǤ˵nm��-@K;�-�L0�$G"~����j�3{�Ke�7����p1��6�ak�Ḹz8�������3V��t���wG�ce�����_.�!�"�(�6A>�NUAg)�&n����远��|�Ɉ���mĶ���:Q����ը�N�䏵U�\Y�wذ�[܂�yE�g��Q��{�J��Va�-�����Qm��E<ُ��F���'�AV���������Ϡ�o�c�%Y���b������&l8������ݣ�c~�\�����l�VfcAi<U��&�����F�^�@�K�I���A\k���$)ͨz����`m#V��C�L\XZ^'�a�
`�)Ob�F�W�`�7^��`��6����jJ��da�}o�FM�J��	0 �ED���������9�n�ؘ�~��v�ۀ�t73�A�?�k�s���	�wC�,�e�1oy�~hi�]��!cXu�0�B
�"HX�S�e��1�YC�3�X;.��&̈́U�O��#�Q	2\��U�5�E9^�~�>�H&�_��9��6s�E��fE�
��P�*;��v�u�+.�P�����~X��}J�B`��JH�l�>*��Egb�[�s�8�Z
iA����q�o	�t]9�0����[�o�?���������\�}�y���-z�����~���~�PO �,=K&�`��>=�;l\t}�������j�+q	,q��ݰ�����dP[��l�6{]*x��I� �,��Fap\b��P&YT\����ѴՑ��K���sNJ>]4�A ���H���K'g��/��`ws�M�s$)xgY~��i!i q0��n |��c�������G�f��k�A
ʿ���>K��E�p����X�b�M��P��q߽8*�=[����,�������T�4,W�e���D�TiV� EU�F'��jmm�SM$���`�l8�ĺ�ں(����ֶ5f/��'ӈ� �^	���0�rb����E�T¹�ҙ�A�i��������lcvsv�E{�5�(hn�:���i|l��বQZ�>s�zr����?6�pey]�BZ�4S����$ezG7�_�^��m�6P�T��@�zd��ٚaER�"��U"B���aoje�� y�G�w�ω;=\���A�)�9b/\��Z6��X��e�<�����0Wz��-�]Γ$�P^j�.�VXʤN�o���p-�}PT�0��Z R����*0�5�L��ƻ�����A
�1)��T���k`�x}�^���:��?�lj��)�)�c��31�̋~��B�M^Uc49�}(��j�3���^Bh.�O�%��z
�
�f:�S>->G 8���.y�΋�>	ǿ�w0�]F��Q�$��-��r$mںk4�rp�r!z�=P���pŗ|�+�%��5b� rC�d-�$#
�mΌ�����/�f���9cߙ�C䷱!+(�Ge0h�BD6�F��k�� ���=K��N?x#�5L�.9�,�M�X�tխ�x	����$m���>X���&ud���~��"(5���Q����|?����툴r~�9Nu�a�|
����¥D�� -2�Zo��+Le�ܓHKrB�x�������4ۄRF��"C�oIֶ��\}���K��dB����h{xw��T�gM9��I;ӫw����Xqs���*|�����}YnX65�#����)����g��G�����5�+���鏶9O� E���a}d�X�sY6	�q�&�K1��1d[���<���u���:%\��߄�_+�?>�|���>%>� k�<U�b%Z�&W�������#3!5�UC���̋h~���q�>pf��x�pn?��ㅬ~���F���b�k�����\۶���5�	��Z�,����{[�m��8�K�HCzf.ѧ��	� h ��f�0�W[�,��f�2}s_P�0��Rs���P};C�UˋC:A�z�cb�ѧñ�6X�8��~������B��o5����c~Fp��,��'����g��T:��Ci�N�G�K�.��M�+�uy�)�:W/���n�kً��j<�A�P�#]0T:��ܦa�4> ���D�-��@]���Z����hZ���y�VZ�^��N�q[Tx3)9���<��`'��n}��daRP���੐����M�V�m���!��s���?��;�VA��\m�:6W)RU���"g�)�p�&�j�N^I�O�+�<��.�S���fM#�d�H���ڕy���4��v� :�F��$]J�	hQ��k�O��¨��j�)s)O8��PS���t�4.Ŧ�>�ҿW�!���Ũ��"oP��S�w�k'=$��R!��2/fM�?�} �P�9u��6�HCj�"�R9*DT����kW3�o�Y�G�Ea6�
��9��K�^K�{� �/p�����'p	Sd�@I�M���[�����~K �$�����+5W���-�;�o0���=�3X��)�l�-۶4��TF��i=�X�������N��{�y�9��H�<*Fy��H����<*nz)%�{�7�1hGц�i�s��TWz��4�s���;�ʫ|��E�
�46�<ydі�Ep�����R�h6d��}^u�ף.�*��N�T~�ѣ������]��m8�\{|J
���LX�4p/Ǵ�8��~�߻¿z�sȹ�����i�u�O��~�I���A_1P�lE�H��<��	'�X���rq.�Ճu.m�U1uc������a�Aۯ@�w"v��/�*�1�7�v~Ι�p�����r4�f#��k�}�W�D%T�F����&IZ�w#憖��hs�1�^��x�氁��t�X�,�W��B��Us\����k�D굸�(�����V��#�+�ȴ��~/M��抻h�G�f��@�����M�"g���!̮uP���Ԁ���V���Q����
�o�zDɃt$�Q�F��>I���$~~����������<�#�tz���kkE�u{~��j��ƓC�Ѯ��"�����x�	XK��	��S�w�ӊ�6����$~-0D|ݙKdMĭsS�+��,77y����aM4�A�i����,Ib�⋤ZR�U}S6����E��hݭ?_���
���d�9q,qP��I��2���P�+���FQ�;�Lp���Y<�0Z��_)h�58�&�s�,�P���rb��H�z|�������a�������x./R-I>�
lRA%}����K�/�1��?�X>�`
;�4��K$s��.ip���
�#�B
]�3A5������ %�W/�-����"jl��P�i\�j�߭���m�j��Q�m�9*J��c_�O�:�*pz�d�$ӵU�8�C�H��;�T�����+�Z�B��0e�_󕨏�;��\�-ز-�&�����N'0�Z�)�Ϩ��t?�O��,�[k�MUϫ\>{�7�dK��G�GwlJ����a~b��_6@lE�&}�������k�+X��]��hdГǼB��26���jQw������
�j�E��|3`4aC��І��b�lEB��̘,��br�(l�;eW7m:pG��Pj��0��I�-tE+��e2�B����Fi����"�Y/}S=���#��@,͕���@*(�ȿ�X�R���*���F�ƨ�o�WO���>�+�d�����CS8�3�*���Ï���Ȕ���:�L����K�ߣCc��k�-k��\ rǡ�$�0�j?���njJd\@93��?����9��bl�t!�f*�Z��D��9<�{P����9�v��<i�{�8ާWi�2H9����0혊,�-�ؒZ��� ��m�>�烉��d4����݌DԙY�p��+�*�Ga(��$��6U��u����y�zԱ���y���j���{.��Z�FH��(�P�O�����ڠ�$ ��B��x�ͳw����4��T�w�
&��T��0l�5jٳ���r�.�L��SQ�񒔞�ά�3�4v��5��P|����t�!��k��y
��{g4C�F@Z��S�m�Z��?���*�O�t�)����x�Գ�-�A2`4[͛L"��B�k��xf�ы;9 �%"�� �P�@@:��^����B�F+�2�fNP�^�2����8[ؾ8�;T^�A�	��?��n����vԯ�����m�E(�*�
�i�m��Ysf8�P�rL
ʩ��/-2zsRC��~�N9�� �Q� �{9�-B�!?���EY��.5�N'�>t�N�#B���[T~�Nܞ	d���ي'��	c
׷�����s����gH��d�N<"��4���J��¸3�!��'�p���:�ꋮ�P�̵����THxEAC\��������ȑV��[V��*��}E
h�bzT��r��M���q�g]\mSZ{�\�لɍ8�y��f��{�Ϝ�w���t�Zk\w��������ErK���}Ah���!�A��a�Z(�`d�a�y�@BǾ�Z<�T�L��I�"���v�j�)6�
�}{3�tD�D\��Ѫ��	q���|\�c��vT�I����f��aA��k!������z���_�^q�`2�F/�>�~�[�va�O�c��B kRh�0r|�.ݘj�N����E$�@�x䤓����ܜK��F���70'#��qK*�Q�_�L�_�5���K ��?��>w��d,�t$3�!�}�N��jo1��2��6�
�g����R�+1o��;���(X�P��SW3�͢9Û����}Yb�����x��P���4��1�e��`SS�f&�v�I�wv�܁M+i��h0���Tn��iE�\2�,��M?��l.D(7#�א<����&ֲ�b0�@Ui������ �ze�	L@L�ϒ�6�����T�ђH݁�P0r����湰|>A3o���`"��W��<�]Ұ�]l�Æ/O���|h��#nΪ���mZ�B�b�ts�3l�ƍ�/_;�(��o0Fp�;� ��	�)h���S��ݪ��+>��f�s���s��x��ç]r��O��\[��1g�֍z�{(�@�����~8)�x�J8�
Ԛ�[�0�ȣ�N6XV�'ߴ����qU����8�	Cn��Oss� -���=�8U�NhL��N�1mJJ8W�0�h��V�M6�@D�2��Fh��4�ɣSWA��S��N�����9�f�\L��Y$�YҊ��NB$�f��N+�}�)ņ��v����Yd5�=�O���M���e�Y��ZK��[;��Z���g��k����X����H��'���d@��.������F�)Pv���O/�Gg�mЂ���@���n�`�p\rs��$�J�������ײHP��o��Z��Yee�-I��1�[�6��c�)�]5�ao:��H�t�ȱ��߶�2�l�$K� T]<�/N��AT4����B�NJ��\cTCd?��X��Q��v��#�:��ӒH��n�͎���'O�#a��4���B=�]�`>�������ݨ1E`G��q�w.<��Y���Z��^��Ry
W�֕���oӄ�5��.<\��Ei��S�D�.�,�Gq�c�P����\�x�R�#"Hik�g��,)��\���>F�#�E�<�9r�q�.���yd�9�׫؋g~}V�r�/R�go�y��%��볍d�}q0b�hrGZe�[�9�I{�vH�V���B��pIXnʒ'�
�dyÉܛ�ڏhY�oT@�V�p]�!y�XV�����6��ίS�U+j�u6�B�Ξ!Ga�b�ex"K�0T$���(5��
��Az���ɝ������6<l"�?3���=%1���@�G�Bb�M�J�����lD��-�+d�.@�Qi�$<q� �a_5�|��F��ؽ����(y-0�H���;�G����J�rhwa�-Z�3{����Ѳ��[��}��]�(����ް�P���Vf��>Ο�X�C��y�!ވԸ���ܟ~���mf�Rb�}#aG��ES$���@�k�fݼ�����&7qy�A#L�4��HԌ�9��n���B"j�-�$RmJ[ �#׶�a,Hl��G�LfT�@�om�J�?�d�\��D������
* #9���!Of!����u<_��<����|��c-n�ب�.����Ǘ:8V��C�?o/=�׉�%,���F�)V���I_�4^_3q�(!x:ak@�D$�)����d�ћ�~5p�D{c�2�$"!��rBy�A,�rC��j��� $��}�m"�Fɸ�F�M��=~������M��X�掓N���*�༜D�k��r����,'�#��*ރ��褲�ϒ�c����^J[ǭ��;S��GqΉ�T�f��������Ǧ
\� �V����=H���۟o����x`���1�]�k?�H?�����"7F��� 	O5�fĚ� F��S��_�\(��CŸ�(�|Xgyv�(�t~�%��D�eџo�=�YQk��c頕O[⩩x��_�uT�(����7�U�&�B_%�ܷ׺��z�Q��ߨ�'z���W�B�{���p�
���P�ʝ}w+�f�9Rݾ�p��HH����Cy�>K����̌uD�q��r;�d�Uw|����r�%>��Qa�K"s6z=ƺܝ�`�v�<�� �{F��Y��L��oN��e���5���^b�����+13+��Q9s/����Nn��.�L߮I2_[(5�z�3$�<��:��ZmϢL�Cz�#}z�͸�ȍ��3�ق~l���k��k�H��~�!5�*�?��LU;�;2��~W�鐓'n�N_]���5��v".y��"Yi��@N|0=��^�E��$�2e�=��g�q�c��{� A[�X�d0]%b�B��6[���<�G���x�r��G�gp�h���JǖB��J��+k��Z�AÇ�1c���!��V/>f����ӣ��+j$��+�qi
�8��x��,�O�L��jL;����#`�U+�}6�(l]�a2�� -3+��E��7i�����XS(jw��VcOx2��ƈ�(X	H}����!�^�.5N���{£V�"��M��p	M���!5ĸ5���?,�Y�sl�>��)�(���I�ذ��Qϥwt_���}�䰊ôxXU1�G��bv�I��.)��(��kIf���z@ h�Ԣ�H[Un�<*�;�S�:?��� ��%�cVSH謋�+���^�_i��|!�W��YL&K�R��*��������y�i���K�D�����[5�rQ\��+�"��a�v������TM�+<>�8��5o>�tWEs%�*����Sq �9���<LL�	��;I���&��F�߈r��^]`�7��w*�^LO7/��D�'���Dr~��V�޻q�
�Ϻ}�]��vo�W�W�=��o-�z�b�F�*�:4erɄHf#�\ˋ4@�%LOmP���1R�2K�d�)G������5�v̒O�F�w����u�T�G^K-�a��r)����h�X��J���v����#�}"�X�������� -y���E�&W%AM���<�W���j�{s,C�E�V0~��|y�4BS=L��-�f&�j�JEd���z�(�{nJ�<P��/N�=�I��4���J���Z�m�x^ܭRIZ�-�ǘ*XGp=K[��Իq,��d��W: ��
ﮯa.��L��~�wgr��BYP�������(Zzc���E[��b3vɦW�9+�R]Ӯ.1����Йa.�M���	�����8�5'G�&,��S �c�Q�=b�Yg��;���]�a��*��$&c�`�'*#I(��+�٨(�1:�&_��w����~º5x�@��x�:�c��q�[�\�f�W��j@lRmoI.+?�c�m��d�I����g�I�]w<���o���������" ���O�^5گr'͟gcN��Ng�� ��#�+���A>�w�f���Z#�5n*�{(x��S�;��vL�ɢX�ꃨ��DR��)շ��]�J?-����푖�p:�0?i�zp7u��00� �{��ۓ��4�OO;��>������k���b֛!��d|R}�́6�a x?Nw���P>����M��r�r���).|�-��с��bP��>��E�pq?��������ev,V1V)�"LA^�T3��LT�.&ȏ[Y\t���͝8��oj�#_���dp3*&�ؔ��(yn\}��!Jk��.�"��#�Z�3;[�o-^����O���W�oi��M~[��D���� št(.��5Z����ԱKX{)��r$����M(����V`�zz&nG��<����W%��{ǈ�	.��}���1�L����_�q���K
�Z
8��j��j|��Э��Q��̓�ށrKΊ>Đ7h�x��b���T�Z��RD^�`}�HD�{Ye���keg���Nb���x؆p'�(��
�+��CNt�<ǹo�V�T���p�l�\�� a=�ځ�ݼKMG��4��T��O�f�v5�O��xúf�7�&F�(\V���6F\�H��A}5���9���Ą�\��9���t#o�8������PύTz�(E��2��Ī���+�\��*(/{"hLd�>�@�i�Ez�r������&�h(��G�2�]SXd�f<7EBc᳈*�zc�ӥ ��e�fmu6��iKF8g
.��<�����m6��k�H%�2���yK
%���de���1¼�!v"�6]�K7jG	z���/��-��?��"�X�}�Շ��!<���ͪ���ͽь��
�+��T�<�3�--]�$���y,�}/ա��-D+|�kz���p�D��Q,ܕ�gd�(�qY7A���sKv���CZ����"S��tc���(�f{�f:���q'v�9t^���Ufތ�V���$%�{�u����,P-~t�������3(�m3ͥ���|@�7\/c�K]џ���z�4%�{�� #m�Sd�s�Q\g�����/�jC�:�?�٤��$YK0�*lG&"��ALf�����!I`�\�ɪ��.|�qrU��'��O��grϙI��I%�PYu0�l�ʞ�㋸��CJ�Ʊ{��������ysp��`igWtM$2*�!���D�4ȄA�Z�t�Q�����Vkr�qܚ��;e��C��6p����u�6 � ω����}��yբJT�$a���7�K�P��N�kT�P$P��	�������,s���CC=�i\{�F�Mη�1PC��^�/�;�S�(n)��B�������c6P�QSx�ETW�iʾ#:�PIy�6~{���tc��D`�/����Nz��~�{����VM���TW��롓"����!�N�fY�5����c�{����;*&_ qFoR�h&}/U�ū�=�N�'kY�D�ܯi���P�0
�/�n�f�	?jE�D��=�0������4�8��[�P�xP��Xr�(�:�X`�O+pF�o+����)��Am���R#����y�P!%�E���~���������Qd��h=����0BGUg���j�cĀ���6聊��{i��p��V)���iE����XlʒC�����h&`�#'NM��N}�_ȥ=L7����0q��S���>��}K!����e��4�4���ߴ0��E(~�/(q�ـ����{v�c���An5�n�2�C�ێ�D'�'s��`F��Nb��mcO�S3�xyV����,�e2!_H �)Gv�����_���踸��=�U��DF���#�1pS�$B#!'e6��k�C+����D����o�')7.��Hq�A�d���Xҕ�[�9��4x.�y���z��tr�s�Zgr����L�ƈ�7�&ų�(��0
��}����L�K����f)�#'!�5ڧ�e�c����v��L-g�<2)߸o�
׎��3�?Ne��l�3 ��,��h���� ,��QmA��t���O%��4�R�/���������،�(���7���|6�%e����s$l8U��yvy݆=6B�F�:)hU�A8(�-�R�^�P+H�f)�9�CG�ea#�%p����AS�ԶN�������d��4�O;����� R�>�zM���:��5xg!~a��k��}��F�N���#M��VJ���12�:S2�۠��r�ge�)A�+�2�i�GG�4L�.$�?�L�}i�̢UW������'��4�x.+L�W�:]{�Se[�uwg����i�'u��Z�3&P`lJ ��/�0����>	I�h�-�B:T��De�����UhQ�$�>�V�w��%N�^��2�S��	�_�y1r��^�O�l�j��竏ƮL"��v��S�_u����C-,0{	��ue�:�)��9�i�q.��I�p�]'5tp]v���g%s�*��d!�iem�2K��Gi������9wnA/|d'��)���Au/���&���7�����oueA�:���{�|��Tv̖������h}^1�bϮإ����Xt.��U2v�\K�[�a>�F@i���F7�%��f��������x�zt��Q�G6;�Qi�2gM��茯�d��=m;�����>@��8$n���2���\��M��Xm�&��F�$��M	��#8%�3
�d��d�NQ9^�zQ!X}�2�f�f?��3zgu�?�.����#���K���]���-/s�K�I�j�Z�^P��dg������rcÍ>��/?!�r��.����s����l��$���cz�T���2�%P*o�zk�|p�ҕ�C묈WgO���p�Tq,_� ^�R�Qh�x�U�����vע�a6�r���f^3U��RfO�Y���`�����|�;ٗ���1|�eS���j:+��r#�����`��M_������R������ޭ���9L�8̽{F�sQ�[�/����ӊH	�����d\oO�RM��	G���wªA�}^/W�2;�N�������L17�E��.L��j�/f�)��^����h�U�ܛ�/f�ڼ �R�"n#�C��֤[��ب�'T�������ґf��v��w�!I��x�3�VK�#�{1��;�{��s��Ua�՟���� i�7��}v(h��{��dW,U�!�cu��^cVA����D�Ʌ���ˆq�o��`s�Ӹ*R�����B+#�"�|�����]���~�<\��&��CH꓏	:	��H�,2+e߳�4*�?��ScI��ܰ��P���6kY%e��kVlOnH?���F���G$=�z��ЀC2����Fp`�: HU����N||1e�p�7�B$���x:;_�p�}�R�M [�2���c�8�j@�,�����N���L���?{�'���v:�?��S%x��[g�
Dޙ{Ǒ��Tq������/2�!UӨ�nzŀ}��k�,�K/�~�W��6jrU�Z�pB��B�x�1y��T�+91�m�5��ֽ�V�B�+�x����yׁ�%w�>��N 
�Z�u��Z�T.�ݜ�â�}|<�i:9�Ι:~�Z��UO�t��E��]d�#|d��MK���'�r��9��n��s�?�W�ܐ%��!�%�%3P��������Xˍ5 t�|��9 ;o6,�E����\�4q���s�\d-$_�'tG�2�}oss��.,���R��ũ�Gɘ����9��;�T�`����c��l�~sa{!�������k1��#ߕ��Q��wUР��m����1N����ĳ���jc��2�ȼz���x��2�q�~�?��O�ez�o�н�ʻԯ�?3z;=�Ԫ��V���D���2_��'����E��'̌��#2��&��kf<0٪���X|�{Iv��.}��U�j������08��������3��V�D��a����%U ٢�;.�v�:`>�ah1,b�W#j����S0)��_�cN�8xxSD�3�KT�qsNI	&T�wy��!⩭^$7�N,�y�s�Τ�����+��+B#�ΠX4q뒼��҄�ʁ�ml�:�5��u�����٧=sW�L�S���P?�m�H��E�����1���o<dvA��%�q��Q�!�蕭k^O�%$yTU����
�s����$9cEn��UD��������$�Or�(����څr�Ғq�Zu�
����\o��Aa��|&-�>�.-�[ʹ��z�1�K �edU9�r��ܔV�N'eG@t$�j#��n�o�"���!���zsNN'I�����O+��0?��@��e�D���,>�N�FŪȑdq;n�f�M���M�
ڛ�{Vqn�3� �N�/�ɻA�u���(�e�m�����<q�S8��PJ�����\��������&(A��/�|�4�r���b=���*����Y��iNP�ī(�������@����[�@m�.!��Y�'��.�lӉqň#�e���GÿK���Hm����+�D��Z�̉�B�U�gwC��xٜ�"+����-��� ���$
�.b㻒���ka����AB���v�����n�ʇ؆[���|�*���!謼�k�I�eu��E6 ��'����^�D�'�*��a�ȨD���`�L%��R�RAꦆT6
�n�7��/.��ϐ<ce�t*��o��qLu!x���`PRR��7�U�G��=Y��xDf]W�،���Wp뻔?�
Qs�I�(0�aÌ���7��p۬qfeKp�������g�MC
ƍ��y�W���Y!w�����ֲ���'6�3��j������I�G��?��� g��zaJj�%�����7^cI�X��U{f�Eu�t�hlG��K����?�Q�NI���1i�`� 1�l̋2�U�4�H������c���ޝAoү�c�L2k9��Ũ��IsP'�����`}RX�فY�}^j��L��q���d����H�6�H��6;ג�-��s��6��ɀV��j¥㽹[�(V���TYr`a0�4�E�>��h��S�\W�aG�Ec�.�����m�_φ��|��К���X@�Q��R,:� Ѧ��^�E�\�A5g��Y#�2�b���&�+����
�T�-�W^�+�=b+�G��f�~�R܇�!/�p�YA�ɧ��{�J9З���ދ�L�؋L��{�M"��X���t���Ҝ"�6'~v�4��!��������އ��-���g�N�=`/�2]��p\��&$�}���_�B��*�B#G�of.s��1�k��~y���97�n%�5���V�D����a)_�0����N0�ɯkv�����ڭ�DL���BN�;��潏8�}˘Z����RJħ���L�ִN}�h9^��>���>U��|�`���on������W�5������u&�.��+�ѣH�����(�Q^��]��L����;��Q��ұ�8݃�趉 6����k��.`�*kʌˢ�!ha#��
����k<�"�`~cѬ-z�U�Q�=eE�T�>�T�����<�p��R��`V��s����S��?���妤��?[/<�B�[)srWf�-�=�ֱ�������^�,�W��d�b��9�������6Z6�w?����N�+&�sIV��q~9�&�$'](�f�/��~Go[2;��7ȿق$qh|tp���e���=n"`Q曆��tԇ����BU�7Z=GI�θ4kE1�B9KՑч�<F$R�B�B~�:{2�H֙��z�����j��1�G 8�Ǧ�3��Ƨ�aNU�I�0%��0�a��s�~���\��uHJ�2���mMdb:���5�L_�Oy¯@�fe� ��>6�m��)�2����G2�"7\QfU��3�G��#��t5AS��&	4��C�)rF�������tN]S�S�^��z����p�a�!�EaRc�O�]�"��a~��.�.���ԃ��?�B�K��o]�%09�@5 w��i�y]n�d��Ub��-0�G�&u����_Fr2�ZR�W�;L�p�][�S�@��[O���5���[��!���ɜ|�~��T>����r߇U,�����F��/)
��̈́'Cķ�����oW��gVI���}:��H��2ؾ^m$����Y]ln�Z�ٱ:BAW,I�Ar�˹���d�;�u2w�m�!	�Lg�ȐyD'	���������q�;.W��XX�X�oWϝH���|��a�=�o|�L�D[����F�/��;8��Dýʗ��ى�נ���NHn����V�d�0[��]j��_/2������R}��-��I���, ��OJ0�'�ƜK��_&M=}=[���	 E	���+��v���z1���GϜȟ���V��H�(��m�m����ۇD�w�{s+��:�Q#�����p|n�L���Le(Z.��;�PR�&���ZX�'.+޳!��b�Yy�P����|A8��I���pL���,+���ș��!]���·�+��I��끿���i���a�[e+��O^�vf#�CгG�^��|�U"���3��{��CR�9�9�K�aAC�[��@s������{�:I�-��3��+�l�G8��l�~�Z�W�s�̫4���{��R�<+X�J�n*�x�-J��(g
��OK*�2c���-#Pn�FqL�8'IV�*y���V��`���"�4�QZi��w��t� j1���?�����-&�J��	��Z���������	G�������d�D�I�rP"p  J�d�섪�3��:$|kr��#�p���qOR���(���s�"G�q�Hf�f�+o�)�*�Si���Xx�u�� S,������'w�2��*Ԏ[)�7Jn��8�Q�D~pցq;=8ə��7�~$�G�C�9tK��;A�$,olʗA��~���"]��곡�E��w&0T�����ɽ-��Rl�M��C&;���{*�	`��]/Q �{�rԧ($�͏ ����H���Jp����"�QՐ�]��އ	xѢ������$ `��������=�Ǥ��eC&����
s6_���a�wH	c0!��\œ�v� +"�8�p�GP4?�~��b���7x��~�v�cu>ٮ��K����L�������P4���O���[G�z��~��(�L���B�� >Ա����k��n=��~ŭҟ�TT�G`}�s[?k�7R���X���	�CR���i�ޓeH��HV�'xq�$�(H��0��|����~5N �I���v��sWl�_c9��;��k[�f��"c~� -f��*un*�܎�T/#hm�0�
��(��D����\֬^�Z���)��Y��._�X7?B]��<���~�A�EFŕu����y sd}08p���]h{�h�p0gV�"�ۼ�x/D*�o	�SA`��V(� O�!Ck�$K�O�/dvs��5��������(��KH=��cֶE ǥZL���#I KS�|O�Ϭ��ECc���ϋ�\4N�,c/h�{th_�����(I�G��`�)��x���ܫ��*��	S��b5�g��Py�������������0�2�*$1}�Y�M�w��6�W�	��=z <����t�qͪ${kp:C0���1Q��i��RP���CbSĈ�p���p���}C�<r��|�(����U�j-�wǓ�=��]P%Ȯ�ټ��0�)3L�UeRV�_�w��n�7&aߌX\��v��g��LZBQGr�,��h<��N#C'�Goa+67Up�>���\�0���ϰ1`q\"74p@h��Q�� 0Pa�Ir�#қ>?9	S*��!���8�D��|غ53ՊZ���A�>�H"@s���/�ǈ.eX��h�(������(J��� ���b�XG��U�\�i�~��%b5)�8�Xr.,#��_�r���(3&s9mFa����4���M3!�/s�Ġ��|�Zb�?��R�`$��^�p&=�s
g��,6	+	#�־����®!�k�ASiJ	���h��g��( �L���ց%��f�������1���P1�*��R�xbM�d�f�E�;���C*��d���Z����I�n[�q�a�� H�**Y��͡��b�y(����,�U<���h�����4��L�� r�F�8ه9�� ČÒ֍~���\4h8�7�a� �sΔ�Ő����ސ��b݄P�^�z�G��+Z��$)
�Z��-��^��R����0�O��� ��|�a�8z	������k�O����Q�
Z)o�`ZJ�`�I���c����kQ-��uw �3�?tpjSⶳǄ[ ���{t][�|�Ջ�L���IPX/0vs����Ws���;�x�Z&�K��Y�8�nC.�o`zG �̿������l���DW&�Ǎ4�o����go�)I�l[�q��~��E�������V�.���A ����Ԟ��_�>�w���C��R=����y��_��R��@���^��:y� oR�>�����BDǯ��U�*���?}ܑ=$Js��c5�Fr�'��&X�,��Ul�<�a^�5,���w�>����нL�KT�K}E�?���#^�iE��i�]s���_ˬ��?�<�¸�m�L ��ps�m>�0O�mE���zN�熚x]�Y#&	�l�Fv�j������g/mW6�c-���p2
��$��8v5��r+Ug�bg �h�M����Y�[��5���W���t��� Z� �)d.�?�����ѢȈ_����Eh���ϯh��y1�po���� �w�Ts�e\��:Nd}��[�1�ܒO�����GD��sj�$� -��.J�"���,)��2����W81�;�,3�n���.���랩{T �9�+���Km믗]6ږ$�*@�m���k�������k��
i��BÏ�6��w��1)΂E�ܰ��FNM�A�o/��ޟʯg�MA=�V�ሁN�4ad�n�������A���$�4uڻS���j5��HF�$ �%�r�)�~��lu��!-�j�Eq��a����L�=�͍3�x���?���C������{xV��n�evfU
��r�k�}'O�T�"<9@g��;�
��B���N3~E܇9؎��P2�.��_� Y}�X�V�X��H���oڊHk���`�[��^K�FDGӾa4����z�)�V�
���h�D����࿆�V%�Q�>2J���P~����y₌��������5r=��ӁI��!K����1R^|�6�'6hP��El/��S{~�B���G�TUW:7&g����3 t�M)�o�k�r�%�jCy�+���x��{VO<�b�y(�
�N���M5����X�߃�^k�e�9���:���
�(3��k
t��z����:�V��*�^��\a0�ݤp��tn*��ZJ���~�x�C�`��«�@W�T}�Hq��}.��&��C�۠�(�$�>��%F�m�����d��GM�>b�)�οSN�ր�i�� ���z���mnoP{�N�%��o�t�{=@{\�Mu�Y��x���\/3��b����@�]Q�h`�:��޳%T�k�B�������׀�u	�����+��踰g�;�[%?�����>8{�9�m��K"x&=��aB	+�v�+1����AJa;ޞ?h�l"l���Q���d�bD�� M������61�7CE��T&�����~|�,i�ҹ��f]����@i�t�/�f6q	7j��G�8ϛg.��3cgNG����[���K
]As#���y�/\
�W ����1;�kU�Bx���T�f{{\�:�;��U�T�-���|���R�����;�b�\��H� 1'�EP��.��.����ݨ�]��:6���4yKP�8~����A'g��I��Aڦҩ�v�efv�$�y��|��g(�D:DM��y�y)�|/�
��o��w� �D*�Ɗ�Sx��.+G�ݙ��h�hh�I7�}�"�ʸ3��Ze�]�/����y���`�6�ޯK��:��+u=M�.�8������0�hJR�u���$�7���2qUN僶x�,'<����2��]�/���8�\�7��H�mq�|�'�� f�����0I���6� ����v�����\�e~܉�H7f�x����I�!����"��X+���J-����Y�>���%�*}��nL�	<s���Ut�4��9�����e@'>gX�NI�N��?vT�U�t�g��$
-D�%�7T
�s�t,�Ȁ�cU��#��/���p�5�;g�A0!�sb,�Մ�K�4a��e/��U2�x�}�K�� �OhH�.^��:y�I����A��`v� sr�㧱�g�Lf�_�%x��55(3��P� \6i~/kg���7�;F�瀬��\��:˅ף��hy�;�/�z��Ϩ�}Eֻ��������F���������apb{�|�{� ��M��C=H�֋��?-�6����& ��{����?q�fKK��HnI}��Rrb-�2S0��3y�H���_�$xr���ʿib��4�k�z�H>���Q1Y�/�S�F�K����}T1W�%�}0ʼ��O��~�C�`��I��Z��Քy]���"E#*���Gt�wqiT�J�J�Z:Kx����յ����[C�pQal��=��
��v�}���_�3ģ��.�Q�`�B��g��;�t�c�r�l�w�P毵�bcՕ�S�'�u���R���'�d�^�j'���{I���s5$V��o��~��o�FK�+a�@
H�҄R��J���j_�t�\>西�����o�b��Z���C� �e�SW����J|�G�*{��D��qk��)���0�x�="�Ҷ�SC�]��_���dP��Ⱦ��aL	zF�'ʟ��)����f�ȣ�ό
T�Jg����tq0����s��iK�YM^����A�*}_&K
�d��>E����֡�3�d��м�4᱖or���OTO�􉲨���O ���|p������%����LECR�q��z�፶�}u�;ѩ�:G���<�h�'�~2�\��SaҰ-x�ا�{e	���3΀�׬�3���}�ZU��4��2�j,��Ƀ9XS�v�IK��Hh�L̮W�4�}�O�RΔ$c�@��/���T�5�7���_]Mk7�jW}�9�~ڧ5w�g�_���"�Xj�(�x�s~���~�E��y[+�*'�)Qp��H��D�I�Q�eB�"�5�KG,��*����|MHk�,v�xh���kŊ�U=x��M���#+�@�,�ItP��h��tɩ�(��Rg�e��z�p�U0g	�4���Ȯ�W3Qa� �˥��W!��c�m�赗jҶ�q&,�XrVr����1��UY�y^�${Jh�Yq|5��J1��?��Դ��X�y0\�ɽE�w��f�WK2�5��َJ>��o� �|��'Bz�t�HȰk���=Ex�N�g���x��YW�
ۺ���c�5L��0���3�X�:�:5HM���S�hm��T�cZ�+�T	O��h|T	�l��O�"�Й&�@�#z��B����rj���������eB,��?ÿy�c�N�Zލz�H�7}��� �y?���A��U!y;+e��m�2�F �G�c�/h��T��Zz�k\�������g[������گI�9x�τ����N����;���eH,i)ht�y���ŰaN�C�S�)�/����+Oa�,���ᛐ��w��:I��P�ڽ"�a��@�T��L"��Y;*�CsTj���u鰊�d-m�>D.I��'��W�ճ�N2����(I1]���S-�><�u�ݢM����7x������C�?�������&���c{���ύH��U+JM��}���V��t���Wn՝�)D�t��e�k�Uy���niu��B�o,G�gKJH�g��%�h���2o�A��{p�P��|C㖞[��� �>��
VE��+���КX�`�B�E�O�����m��ݝ=����HC	�j���G@SO�V�����&*�u8�v`��,���t�법�INT�-��D��E�u� ���N�t��D���9�8���y��|��#��+ί�W =��y��@�f yN#��r�El�&({d9|P��7�s�3)|3J\o�k��xR�#��aOvL��A��K��f��?�V�D/�E����W��U-YS	�to�+�@6x���'�ڋ>�;٥V*�H��B�:�)��jΜ�9%�b�K�&5�̌!,�t�o}c+���>1�!w���Q�<	bc�rS��M�� ?��\1*[���1���a�_������,�+���!����e��~�	�`�Xu��0q�v./�� �+�������0��b ����')�����������%5�D����u��"�d�	�C�w����E�C��rYB�3#}._�0��I��J��;��o�j
��&��S߂j�t����΃[.�(j�u�0ϛ>a3�R��ng�m����.��=)�E�̈l�C�,�nbG>1�"�kP~�K��E��xH�VrF
!C�T��t]���~�aP�/���:����<d1�Y�n����ǠOѲ���y2<%�Mx�>ñ��A��l� �q�1"��`*$O����ۿ�ceU��[9�5�ʃJ�6���Æ��r��v�@bI������GVL� �]{�|�!��B[�G�.{�x��@��|V�+��S"|�G4)<������{8|��:�ڢi)%(��MM����V\�xy@�?��d�k�U�t��`��=�Y��i����:A�L˿�Ϲ��I�)��
�G/����h��C�\\
�jm�@��n	��b39�%͗Dk�r�������in�!����R�����x�f<�ѶT��P���<J���ե�D��M�E�1~����8ΐ��_ώ�,f��6\��Ga��N�	�G��#pŀV���N�ۼ�8�Z�b�cH��#l���..�ڻ?��0������9�F�Q_ʄ��j�_-�1�&C?���h��$ >'6U>F������0�P��A��u���ñ�!�y�G4(B>��d���'�@f^��'�tS�7B�!��m|�Wgˈ_�F�O9�j��¸�O�d��6&g���hp-
�	k�@��C���R�5��Wi)=Ч��COz��*]��#{����;�m�FI��}z�1kώ�/�k�� �q�޹���h �	u��ֽb��n<�ƪ#���%;� �y2\W})��`�S|.��E��s'��|_=�b�xE����9�l�
�6v )���N0�f��#���hB��p.�j�r.	�X޵Kk��u�����p��C��B�����(�zNл����h�į'�(���-��>;�M�/M�h���_��P��2� �Vɝj[��_a�5�g�JMk�	�����,�gP����N}vO��o�I�?\f��=y;���JGR�8Y �n��a�-���ٍ���yt,{�r.�.S9U^O���4D�$��ح�npذ���X�YR�l#�s��g!'���A��f���-ZX,Y��N�`�\z򑻑i�!��q6܎��m��Bi9Q��CxR�>�&AO�]hs��g�9EgG��b�[Ɣ R�:L���)|�p_�z�s<���Ph^>�&�)�ktGh1��t�V~l�=?��?�{a�IO���o����6�};�1m\ӂ�W�*!�=��n���Q�k</���f"�x�^lz�0^	x����g$aGq ;+?�a����J��� '�#ƞn�G���U�7�KB@^��|�\����|�뼑Y ��gz��q��U�����9�_d8diĿ*?�v���@5� �
�d�x��i8�Utp[N�چuC?�&y�I��S>�zڛ��;&/��M 8�r�rM���^-�1�PU�͒�JE��_�듻O�L���ʧ�Ȣ�1�_�>�>��^	��n|:4��G��N�",����6q~�V��k7�y(��co�q���4�R�$�80��0y���ދ�;kj[
:�� �8+ifʎ�U/7�-�Pͥ�sԆ���M��!���Rc�h6�U����1Ӷw+���k�}�Щ�hX��u���[�;�"$ę�+��I��.7�ҭ�G�}�Okޘ0�:��x������[��i�νǛa�=���8,O�yx/a�o��+V��{�����)f�MLr�*�pb}+ b��@���m�C]�V����G�Q18������ <p$A�h�.�,nBj����H9�x�i���
�rBd]�C�,1C�P�	ګ���O��zQ�.����î}��,ޚxUy0P�zyw�PI���4\[G��*=<c^�%�`�x>�ƣ��j���Ά�q���ˡ�<J�J�}_Q\�D1r�E�P��R�@��	W�Ƿ�m�M-�%�3�M�7F�ҨK�@��$�88�U켊3עp#�P��o�!ҏ�{b�Xa�|��h���E�� ��N$�1�W,G�Uy�]�f�䧖	�3j��l�\��m��-HOA��У4��Cľ�b��l��$��0�D.�D�ۧPv$m��h?8�����_���춇߆]�)��eʁN�^!�4j�0��<O�p�W0"o�Ì�9\7l�KَP&��g�v����i�xa�!��W����_F�Y�k��n�>��4��
p�Ɣ5�^q�Uy�����"J�zQQ�QUb0b\m4N7�j�R:R91tq��P�� ��h�ʓ>��WaHM��
]�������8�[�$���������Ԋhk7>����	�R�U���C"aB2T�\P�\7:�Џ��uVaW�`���`�_��y�X��6�Ou4�a����s0�q��/i+��9����5N�����
 |p�x�/5�T���,R�Az$"�>l��"Y����ݻo��̕dm]������3����j∱���\��/c�5C#���{�����֬�V`s�s9�B���m���'?r��/9���|6|4��,l���lsMq!qc=YJX�����#ԡ��<䫺��!�n���R�5���I�)r�d�p�/��+�?��B%�d�e�Z~��q����	d��� ����T� C�"��lC'�ҾL{���H�XΓ��)�e����KP%4� 4���z�dZ��Q��=�Bx�*��[�%r��B�����E.��'e��q��������e���Q˱�R�>[��3��}Nꥡ+�)�^_
"�o�.��; �MH�
X&!�MC��)Iǋ5mdiV�6x�ZDE֥���<]o>��لE7dG����R��w��ṋgP�B�斵�X���R�¡��)��"�M!��~)�q�y�$���ջ�MPY�<�h�\̲)�͉�z�H�rr�c����;�q�Ɨ�2��S�w	/-�#ğ�{(|���f�E��4ns��
|�]�c��O�'��������
kU:@�IͰloެ�V�)�����҈ϞB���X�F]Os6O*�XrTnQ`d�r�0l�����]�]5)$��(ֆ��R�q�;2a�*"fǧ�D�[T0�t�!aGd|�rV���u��>�?*�x[g�i��=�ht�H��f�K����|�<gs�B+�`�<��Q��û�[����WS�Iɩ�7lD�Gb��#+�����~ M��ӏ���=]`���r@�;$U�=I+�#������k��W�w\6�FP�KV��qB�u�P�̆���2.���AZ�5�����Ȍ	�i'�<�q#q	 � v��:� �+�0�~��o�~��ߣ"��s�߇�|�p�=�[�]���5��J,�@�S�� ��o��iF�.P��㫦WF�>�p��^eW�:^3m=CX���Dwu�8��҈F�5I��|����&'��i���G�<8ڪo=�a?M������V6@�6�S�(+�5n��71:ϺO��7h9R�g�+n�d����
6�0���@��c�o�'xΕ6W��b���Q>�"���Z�*���'��Sx�k��@�1���t�6�sS�0t����LO��^F6�\��i�
�#<x�l
[�����-3"�H��Or!+پ�a#���;jy�PWQ�W�L�����2 p��t��s��r��@��Aw��LЍ<�D��ǚ��� %��%��Zl��-��sr�=8g�Sz-��ζ��q���z��9��SJt�fZ�����*�+훜�NĳB��gȳ��7_!�P@~��0�{�3Y�wί �T�u���T�M~�RQ��t���d,���ð_���R���+�M���z�2�&?�P}���O�m���M�����$v���t1��;�M�3-�&񆵽��o��#�tQ�hs��
�-�C��@�Ģ)¹~���{؝����������Jf4ŤO4���Mx3ȸ��O�^:�j�����?9�t1P�`�-�(I�݃�?k�5�ܔ��5��� ��BP0��.oG�0b�bOg�1�՛2����a���LD�����������z�TA$[�*��ٳ���W^
w%���ye��l\��tO�9#�喅�cl��]�[?�!h=@�����|��vD�7/�K;���ӯ�6O�bv��wh�9p.GT�$�ۭ�}	�Q�J`�H_�d��i_�>8�3��8K��ȧ�h����	'�����=[�ڍR�&��VL��-?'��R����o���	�
`j	j�J�P4��e� $
W��n�{k�o�R��5S�rK�����Mܯ��[��!d~W��ˣd���m`�e���,hg�2مu�t��2���Õ�^�k�̠�X&'��X1�ӯ�{�j� �g����h�d�6������BB�2M���%߸p&��.JO������3���ɾ	ς�M%���gd.�4��W�w�q�/]|�mn�.:ߛ�?Z�+^����ژ7.����w��d��rX����� dDW����[�7����VlJ����>���d"�X,���%c�c�z�zfH�		e�o��=_��b���)�΃��j.����W���W��'�;4�YLt�dj�;dj��#a���w�`�?��ڂJ�̂�7R�� HG��O^�'��!G:bF0+�g�C	��L�=v5����!���P&�o� �}��
4�ٴ�T�H��fv�,+�m�D[Ɔ@s(BR������4���aQi�� �C{�Côg\�&��3|٪s��F\���V�+�bU~J��e�L��$?���\� �yǆU�5��e�A����*��԰���Kj]|�Ty�A�]���'
o��99�򄠩H����g7*0��V��E�7���4��r7�����h���rD�%��lG��Nr�x��rxd���mHy�����S`C���T-<�Ve�.�"��i��W�7�5(]�J�nӺ��A�Z���*�Vwx�j0G�����]�b���c�Z,^��27�N�]`=��%���KÔ�@=?��X�1�;�Xh8gC��)��6�W�E7���GTW�ܫ�h9y�S�+V}����US��������N:��}�2�ɳ"����̳�#�c��.��邖�_�����.��x\�Ī�oX
!Ѣ#8�A".gJn����X`�u���iK����H��jԺce+��z�3�eR��O��%� ���џꪔ�W�3-��^�U�����
��%�q$�#R]u�,�v��r��9�w�w3moo�$�G���I� P��*$�}vS�e�O�p��k����u��V��%�ӢUa>^W̋2I��7��xx�q�bl�nT�)p��)�#�4���������طe8�x�@����ݶ�'��Ð9*�@�.Jث�Ƶh1g��fR���X�<����]F��}��M�;�}s*�f�j9�o}K�*�os��]�$�TX�h,�g����Ö�#@:s�0��'2W�x����k)�@���w�ȫ�t­(����`�
1���,1�f�� �H�z��k��Ce��2�|.�����3DjL@�n����t�S�W���3�b��L!��Y��~���Srw
�p�n�]�ywŏ~��7�mh��'�|5�}1c�4mk��0��^Mn����Z0���Kx2j?$��WxX�A�k���h��b��#��?˗��P� {��J>������[e|�b� OȺ:� ���4����������埋b>EMLf��U�\Ȏ�S�2�)���h棬i���>U�g�\��΍�ӑ2
-I�n���Q$E3��w/���?�;�:�?��P������[�#��@��3�6�2��`�U��|���;G���X��-���>dd���ξkw݌Há�G<�P��x�Ԁ �t۱��
[
���Xe�I¥��r+<��/�(�C�
:��Q�݈�#`f7˳q,U��/��0��ɌR��r�gT�� [6��_������tŹ3��!�����`���1��WB���ɘ��.o�_��Õř�P'���h-#!��#VN�5 �]h�W��_���d��-������*�9�p�XLJb< K�0	E �~"ρ���Ӧ���t��F���!op��-�@PK'j	���0�*�Hy`A�@�k� �$�~'�!*��n��V�������� �47�'�鬆왋��xb�.�G,�W�9�=�Fi��T�	��ԫk�儌E��<U/�����P��҆��~!�݄���S�L-P��ʣ�P_�����@�?` z�<�@E��j�.}��M�
ߕ����Z��>��Z��N/�v�+C(��?�����T0p˼.��*S�7��?3����vZ�g4�.��Il-9wŇ��t�����:�G��e����������#�oo���1߬���q'�K�ɌF-�:x�9;�DƮV��C`n�w�/o�m*�^�S(�/=�8�K��%5��Q���\p)�r��.�2�A*����1�Wxk_	��e�T�K��]$����	������f��=n��{���r}��^O/N���I�H���d�KϙNd)�e��i�/�[ ��T��֫p��0ܮ��ka���k.rb�������<���ݴ֫��P�4]h&����,s�<3 ���ȼ���⣞����N᨜	b�Y�K{LYo��*��q��Z�����H�S6��@��������Qp�OY/f��!�S�T���OSy#Yɱ�:ƻ*��w�N.���3�pq��[6ƿ�a���-ϼﻷW����k�6��Oi�xՕ#�$�l�H�0�Ԇ�
�C���9� '����Ƕ�"��%��E�R���}1ib/ʐ$�z�k�!�S���Є�\ �~օ��pC�Oh6%�k�b
��@�Ҭ��Wpv��������io��gq���Z^��ȞBu�^��J�������GgO�#Z4�_hW}f���K�҇����w0�-UNi�H�U`�Yv\E���>���d$��c�>іݠ9Ņ^o��~��1��7s��!��!�f�6��	��8I�vK�AS��:�d������rh��or�w���a/�'?��.}@ �#��_{��,Z��4�(9�U�<5�h
5�O[@���Ϻ�>hEh\<�E���*\�|��!JWryJ�|n wj�>{���kʏU��N��C����SI��^�m�y�O,E�lQ��0��w���9=Ϣh�pD�S�2&��(Ҭ�G�{����[������}��(�`��)%W�������Xv̈́ENԛp�t�NQ��u��nD>c�.���2;�
�bӷ�?�'������n@.��H��=� �N��=�˩Á�3�	����Ok�J-*��DU�
�v>�
�Ta��g�V�<ĩ�j��~wGSH���H�o"��+�rIn���n�L���K��Gnr����Q��Y�3I���7mQ�k��n��x��<��E.���6��H"X;��,��
��z�.B.�q�C������ r �{�:�O�Iׂ�Z)T���ƨ:ˉu�����$�ԣݞ����=��<I��)��˨h��h�D�(;
:;ޤ?��=�:�ev����I��4iaLk�����9�%��6sl2Ey��bz�>�لe��ag\�A�=��Ŵ�v��)�+kƥ���K�MLiMT? %�B���X�a�p�9�,^�!2�l��+�U^I㺅M�b���c[�l0%O��LT�.z�v�"蒝��P\ ���N�%F��g昤v���AJ�KuD�t7`��=i�C�!�����w�b�Q1�L�ֿF� �S}JN� ',�D�**n���s/g��7�%�:�b����,w)�mK9��NϐN\��K��F\&�H��+ ���r����5� sK+O�J**b)\���|�;#nv� a�������՞��K�!I��U�"�wpE~�S���}���bB�?%p��gq5��芬�7a���S!L�b���tc����G�ς;Ocm�o<��������6ɦ�9L<jo9\��ˑeגv�~ٮ
�Ã�K\��k�2�x�����?�Ԕ�ca���xx�Cub��W۸�VH��Y�e������|��S�J���>v!���G.���(�|��r:��L�O����_�У��}�W`c�o��1d!W'LMJ	Z�5�"�o�o*�c��� ��bg#�[�*��E�؇��4>����U�,��>T��d���B�;Q0{���4����0�u��J纚�����2ۣ�E=8��1t*]�m�:'/������&���[���Y���Yc[�\b��D�	��zy������T����f���ʂ��ݟ�$X�͊��c�6ę�Tdǘ���:GYo#�`� �����C��p�JЀۡ�%! �j(l�c:���nuª@)͕�����90
i���DD����K�5�[a(H��U��[��M_��w)��V�ef"��'qkR�/�ɶ�Ȕ]�=uqX�蘛�;.R�.nݤ��9����"������Mo{���^�U5���k݌^ָ,�P'����3k��'�X/��L���ąr�;,�b���y�}N��S��0�4�6��ƴ�9M'k����*v�6�v�}���$���3�X��u&f&W��)�x���%��|�.7���X�Ӂ�Ｉ�a�H��>�3�tV/b-���udKO.�&�0R��PC�qPQ��%�C��k}r�m�s�_� ����:�e0��W�w����ΐ��\Ӡ�o�J��Y��)�qN�穱4�M���-҂?v�X��1��F����B������?M��6LM�7�~PX;�����*�g�f���=��w��h�⨢E�Na���M�}�y��D�iEhtL`��O[�����ܟe��V.�_���aȹ�ݙ�5�!��ܥ�����?�b��X�9z52,)�Əo�`Y���X�a�����C3�+��~�%8���fe��ՄS?��%�`�U�^K��������X�Y(��҃�
Pb�SZ�'(����BZ�R5E�vK:�|C�F���t� Z�.h2A��{a��K�����a:
&v%4�q��#���o��5C:{N]?���o�}7�M��ZJ�S����S�t>�$�.��/G�t�8!H���.�F�XRi��R�!�9x��GC���w�� ��T�~�{^`��O�B��嚼 GPwnw��v�aP�ϒ�W���(4��L���iz_R�r�?F��<�+�M�y�njs֫���Tv�IN���^�sQ�48{!W�gN�q;�e�9���[����~�|&xi�o'q
Rth������l�A���DN��k���a�k[ˮ��R8Ri|��9���ƥ�����'���t���}��X���s*�����E����1.7��Fbs�@~L��,�e
���)�����GB�����RC�5H-��ܺ�BL�Qc¹��r�����s����m�!;� �>}2��"�D�|A�w~0��\�ߤ�S唩��+����^9�\܃�9E �T=���x�h��K� �D�^��4���4"� �Ъ\�^��m�<���:��ۏ�T'g� H3��K��{���X�SY���J�5k��(k�q�/S<�S���+sE���[\�]�DQ�ԅ�@Ya�<�%�j.���E��<����j�=�%̀J��b�R;�rǦZ���_��93dDC��#�6��?���ǃum��`vϣ��Vf�Sq�J���z8|o���ŋQ�e+���NB<l.Ng�Ħ�����/���P[Ie�-�L����~7/��OJ��p�����Wk�UP^�)}��)�2��h! �[���v�߻<݉�?f��`3�i��>���p�L�R�I<�U.E�� Q���~E�`Ǣ$�i���T{�&r�J!|���qm�}*�\`��L�6j��Q�Gf��^��CR٩�^%��m�p���������F�"wj�P"�vىEP���g.�߬�t�1l<Zc��:e^�d<�����[�W�c��1�{'3�˖ib���+8���	�B�~�v�"�/ρ�v�Ŭ�{7q� �9�.�u<��� �2���� �-'���XO�n������A//�7'G@�Fq��g(�C:H ���͊�7�_�ϊ���R�x��8���SJx�|�������/xL\OFwH�C�@�qo�_�f��+�	i��pr�Eߞ
d��3s��~�g3=ڻ�!�r�"�ykm3���W�RK�c�Z��LY�/P���N>��"Np(C"P��=kH
4��8??��0����65m7 �s� �59��U�c�������y15�(é��qÀOԺN����e%��QMk�:���Q���\�)b�i�#���ѣfv�X�Q����aV�ssdx	*OV�J/���_F�|�����6��:�5�U�x��z3~z����e����1�����X*p����f�e6����v F!z�zZ���PAB�X�3�W�f��|=�oKR�N�����Ak��u�z��5��+=��D��g�wg�%��۴�@QT������y�|�֥�E�z�)�$��I��zB��k�U�5��F@{^yC�eq�6�>�\'XG-�1[�P�Z�i ��0�sDօ����r3��xй��K��˚] ��P��È)/���ை��-�I�r�,j)�_��� ���a觜�Q*VӐ�����#�����⩼`��
�M���H���M�u����xH���<����������oކx�z����E�^���B�v?P����;�����_��y c�pX�pm��?��H��RW]��N�j8ı,d}�	vM2�]����Kd�Ҥ��PgIT�q𕢃H���K�������|��?���I�������=1���| ��x(�D�Z{�J4K�O��n�;�	�\&՗R\��H���C�8*�� �������k\P�@'K�bkOOl(�ff�bڊ�1FN�f�І�<;j���/�k}�Ǫ�x��<~`>�'��~��o�UAG�"v������MY��;y�s�1S���%�I����f|K�?!�I��`�m��]�0W�zP��V�/��=�T�O-3��� ��~.��J�Ai�1�ѳȇ��hD�̡��p���:��8�%>�o9e�&1Q�r'aX:�4��_����v<�d�����&y���Ff��ڬ�O�D�(�+����n��$D�M��z��!�p�9������!}*��J�L��>7� ��cNI��s��L���C
�p5'� �����Z��2n�?�uRu��<�00��(W5	��l�/��wy�������EӠ=v%G��A�ӽ+�J�5�\9^&��1���K�pNdvT�r\�>�����y�c A��J9n	`Z�tJ¢���xvo��a�l���?�����NQ��i�Ojo�,D�cYgm(�?t���/#<α�R���&�^)+�u�]@�^2ͳ���V������cM�
�A���O����z;kCL+�<l���Z ov�4�Jf�$��KA��͑��p��k��P�;��K�����!y�KZ���E��fB�P]�}(xU�䉗A�͌����`�p��~�Cz* �FP��9���ChB�E۲�KJV3�֓U� Px��@;��tI��o�u���m#ovb9<j��-��!���g��B&��@ր����=�ﱹ���dS�����]��.�`Y�'�հ����9:���z�q�=9FW���l�����˃��*� L�2 }��0�d��o-Ĺ�>�&�y�.4L�ބ��y�Zq�P��I�7?}aI~K�]{�%����n�8ل 먪��US�ȴ�0�<u��3oq���<
Op�]vf��2y��X5��!8�t�5��ڜ��(Z�8�L�DV$�R�SCix��
6���b�_��%-�:YDG�ꡃK��ٵ�RdCYҬ��
���ڟ��)V,��U�uSD�b_8J����͸�
��/�'ިx�m�#&����]��+���;����Ҏ�ߛ�Y�����
Kot�����25E%r"2߶�����3���m"�� H��˪U�
������>[x�QoAXD�Gn-Ɠ��c��T�ja�P�p	��\Uw�j�9m$��. �Q'b9q�;�s}lѩ3�sF������/���Ah�+��QJDH������1ۣ��B��uj����qUͤo3��j��.�:�G6F/r-�z���σ���}�}�8�C�?=�=����{�9^�:��(�&oj %��
8gIi��ef���B̤�M������ -��]Ad<�������UA�ݚ&��ލB}���$2U���堐0�+#��9 W1Y�r��p�F��/��wD�ɀR�v��̕@����a���;���~f�4��h:tgm�@읆N�7���E=����_3R���yNH��C��<�źD,x��^Թ.Ϡ BW�>W�$�lG���`4xʺH����{���͋�eڶ	L�(�Pti �q���@�">���~%B|��z�wAmƇ�������G�0a+ڡQQn�&�!;�= 4����wd�T�6G���m��$����Q���4�h������{k	�=�-������P}V�����9�'�O,�.�1HC)���L!Z�%H:���:�@^��ʸ���<� m�ʦ8%!��G��T�� ���q�<-�xU$Q�_G��i�Q�39��?5�q(�C�g�Dٽ��<\`wR�s�/f�Fy#��:if��YF�5r&�E��Mm�(���vY���꘼����rr��k�w)��+�s|-B+C�X�At'�`h
w�m��M�6�*B~zg+�qnA�~G������ߒc�D^�w�~�(����S�����eC�)p��k��y�تnM#���>b��.=�Oݟ�x�hd��(���|�� ��}-��ѝ,���h�g�M���t�'�8��FZ3f�~�"�YmĈ�-4�uP�x������V��N��za���Uu�6���L�A�FǳN�2K�΍��-�E�D䰗>��n����j�$e�Qtz�:��Dq�6w{�0����7fE|�.t1Ԁ�%���V��&h��
�e�-�`OWz������4qf�11e,�߅�r)�3У��H���p��'�� U2e��W`?�ߌ��p��SXa	)K�Oa���=�2(S�M43a�ءV@*�䳚�(nP���7��.O�G:��	����Z^9q�Y���[j#�:�s9}�D��DT�I����X�7��޳}�>�n�`xe�j�,���~B�[�����+�dP}4��~���&O�u�1�2"ĳ�y{~�\���j?��..�#�u�CyU����S�a"�y�n��'�;�KՅH\�y�}����n��u&�nX��[�Kf�q�ʠFF��3��&o;�wX�]E�_'�Ҋ�ϰ^�`͡-�7��^�J��K���5�R������D c�Y��*{.��*tΘG���s8
,O+�Sa�%od
�N�����_5~��Dt W��������t��fp���G�c�IN��M�����遇���sz��j�Kxt3��"!�{L�m���]Fh�+��	ޜ��B�����ɍ�A��9��v��gB���0;9��Ѝ����?�s\I�p����<�=�V��~t�� ��4ʳ��_�V!7J�Q����M�l����,/�T��P�S! w�P��:�af�T	�:��NN�)�����)��	+�p�'v�n�]��w��t(RL
l:u��J��Y���Mۢ�x���oz���᪒�u���(y����ZK/�L#b�����ӲT�6>9,�w��Zq���Q&�,YHn����q�2���W�tA�\u��@r����q�(ݹ�o~�{���K���2��a� ĺh��%��o'��7�Vۈc�s��"�����Fn������oiɰ��t"v`����C�� >$ێ@f�i<mM�ٌc7�<�yd C���FIn;�w�����UMv��6�~&z@�[f� �=<�}h@t��ֵI�}֮>�S Rd���Bf�ߓpb�N�i�`�1d-R����0IVk[�_�Nq�al�?�2g�#�?|a�Ī>-'q�^��s�FˋT6N0F��tU�4�U�>�I`ӿ&\���Q�i��L�y`��?.L����	N[lk7�%k�h9~J��X�!7�ے[B?��"�@�eR�Ȫq��`�h*�X����%�Y�+�O�
�vP�:)@����ו\ܗ�p�(�V@�L1��`�tPx`"�{s���Yյ��qU"����br�$&�gq`��!5�1yH�"�F�a�5���i�U�����8�oZ��bN�$iٱK�P���G��n�jY*A�m@/>�4��n�b��
�E+����N��J�=��v[�_r�l~b�F�-�1JG�Wk�.�E٠s}�����3L^LZI���zxy�G�T!D�O�g\nX"BĎ� �YT�;-�e�[Ub��L�2d��1
A�^�M5;
FzY���h�����U� i��b2&QIoܛ����Nm<eG�D�cJS�\R��Tj��|J���Ԛ���1�4����y���ދĘv�+���Z֥����l8Uv�9��m�E��B{�\XGk5Ã�TH�mX:y:���О��y� |�UY�Qܑ��ӌ����2�Зo���>GjE~��M�Cr�A����EʌG��d�_�AAԀv�A������$'#~��8�^�J&�|���*o��������95��R�URA\'���`,x�q������%��2�A������g��/�QlJ%~2���<�e"��g��ɴM(������W;�����`�ì�V����J�p���O������^����i���V
q1j�D�jZ�(�I��Qx��QT�MAX�5iH�� �3.^y(S��韫�g�I\����L�T��wo^~M�9��~��g�q�����c�iM�p"���k,	!�I��a־a!�LB��J���K�̌����rNp���@� �*�z 4呿Էf#EWm�.����zO�͊�m��V�toI�?_i��*qCZ�	��s%(�I_kÏ�K�c��,S �Xo�Jm�V���O�B��I_d����1A��L!P%xe`���u��F+�<�Y��=��Z0���G�ijORD�9��b�f���Y��I�� {~^l�#��D��\�dZwlt���=��X�f��h��9��͞���J%��"߼�H�}���!1R���N~���Z@��>���w4@��}j��6qU��i�ۦ��`�e�7��d�5��zeCtx;@'��nm| k��$��dv����;�<�.C)j(5��l�r[
ܳdH,�<9�c��
���u(ܥ��ɕ�)�?���%9�6>�܌1Ŝmx~5�W�1���TJJb���I�I�ݮ .�mb�q	���Ӑ���2F�"��IY��� D����kyT6����8.eaZ�w;������k˪$�.O�������y+ޕ&o�~�R�c=&�[���8��U 8���3����I*m����Ǵ���F@�H��ĳ0��%o �dE K���%�@�r�{���ٍ�O��Cb�;�N�����SfytV�.m8^ziF����m�@�Y�*"�褋s`�ƞ]J�T�6�F�1���p��R<m�X7sS��b�~�j�9?�Ve�EB�9'a��&!ªB�~�~�=���c��D���_�<��i �v[���E�4(�Z?�h@�zחt^�n�B���3�B���!�5)JT�Q���]8僧�@fb��H�3���v̊�����3Wv`-s)�	�^ʗ�ָR�� ��������/sa�+|bګo�K �*]�MR�D��ȏCo���,o�G�B�v�m��ڞ�с��ow��nD'�n��󎾰��!���A�~u�UU�}���p�?d,Z��'���9B-O��9�ټlQ���QV��]%@Ǉ���U$�߄���ۿ;[T��",��/\�Q��Â?�Gb� iM�*-��aי��<{�}a �
�YZ��J굇%ܘ�g� ��x�����1���_ʅ|~&��j&9aC�Ѷ�.�G9/Y�/�� 9{�7�tn{��N%��U�M�i#=�O��P�D����x�
!�@$72fs|n��6,��,߄Ri�k������R�D_����0���r�-�p�iG"���}
�d2`[�d��B�v;S���"���>��e�f6��k�c�����v#ާ��-� �7��nϹ6���L�`���^�ty��gp!�Lq���ȭP���+��Gd6]c�����=�jǵ�*B"�I���H�E�і��<"�36p�������p�8r�Qը�7��,��l�	H*^��dh�Q�������v�B��l�cvHq�r#�aZQ�a�)�M6��B~��[��&�i'@j^C�C���%F�#�Z���c�:��{�$4Zx=���=�?�9��9%��ӧ6u��0����:S�k��:�Cb(�����+B��H5�s�v�����\Ą/��׎�o����^x��q Y���p���`m�z�P��F��[)���1�,�6?OM�.��������;�A �3��CӊEӹ]���P7���z��ʘ<V����9�E�ڡ�c5��߱��gN��3q��m�t�E;�.��0��X�ۊ�b��aܐZ:�:��co�j�Pm�&��}���1�l@R�1+j	K�������
6��{�����L��5�`lA�"4��pJ�gM ��¬�s��_a�(�Y3����,��L�w"��F�Fwu��B#|{���O��Gr>!��&="��O#�t������#���������D�������O��0/ˉ�5戫?��Zp���qv���t\nt-$�������=OF!b���-�)�����8�s
Og����_pN�Oz)��G����04N���/j����J<t�q������`b�Z^��Ŏ�ʫb��5�LR��9:��2��K�t�Lg��aM$��zt���y������Ў�Ը&?��:�X�B5	��e�O�M,rbs.�8}p-�����`��3��cԉ�ن^�,��|]�-F��Z
{�i��� vS��)wXs��M�X��^L�dMX��$N��$�q�E��)6��4��Gh�u}�H^\�*7�q��T<�Ҟ�\Яrߟ��zY63���c�m4%�͗\}9&@�/���t�sD+2�E�B���l)�v �q7z���s�-��Yv�Qà��ԓ�S�o�<�NP���Q�w�E�(ԁ���=Q|y'��sa�����( D�+�J����k33>�SNt�X3aQ���{�+�M�@T�����nbB��W'!��R�>�.�m�6e�XC�<z�E�H���x�"Qcq=���*�F��fG���`�ޭ�xؑ3��,����%a�΂�:�4[ܢ~���˸�'��S�z���ӌN���_��a�~E�<�1�Sc���,���	��yfi&M�<y�S�$W|'*�]�q�?��Lʻ@��;1t��
�\)�(�$=l~r4zw�w�q�:�z�y@z!�c=ㅻ;�by@����ʠ6����u�B!��g���;�r�Dgm��vzFN�³��ņ �C��*$FICH��ޅ�R��<�}�LC]}��
	�|��a^�(?��G6�q|P��/{�r+�>�%{�U;pL��>��	��V���h"�J�� :(��'�w���K�'�5>K�؛m�\$��F4��>i�#>�Aaּ�;�v@I��v�,'��h�iAj�b�r�������G�}Ϙ}��N���q�~�q�!�3�\B̀�Pa'�/�C�|��~�0�b�V�Em�?��&Ǜ��R%���=�3ZQwOUc���M�w�y���ͣD�D]�_��˪�4��ZL0z��+R�J���nf>ش��0���
r[���{�hW)y��uzw�E��'!�%��J�B� j���d�B��~7E}���{?��Iq���u�"*uO���X�p�'xI��'P� c��y<�7�Np�v��DZb(�AJ(GЯ���?t�H�I��AtDs��Rx���d'l:�e1<N�w�}:xiŰ�� �
�@���8�RM<��"�������T\�Nx�Fǐ�@P�����_��|3X�R����o��Qu��c�L��pJ(��{�jN4]*o�N�1��,J�>��M�B(�����߱�=Y��u+\:
WB����,��W�>b�sC�ýW<J�fK��_B~��T!0X���ѳb��r�*�T!j����]V���`�?ze�������|<D���>r��u(�7rޢx����hCj��IJټ�u�L'����p��D͹�9�U&&�NӴť�sE�^�R`+˔�a�Y�	���ѳJ.�K^p*o ���#�dN���8ub��ꚤ=�W�*�'���3D3�K�v
��>��2���Ō�)��u�X�����@�s�_�MB݉4f4kH#7y#���ϸU@�v����c���G��fA�cl�h[����6zH���;��o5%WF���B��s�!�=LP�ik��: n��
ן����@4*B$ë�ș���w�;F��π.�6�۵ܕ��EQ!��Ыkw	\�c�ş���@zX�G���֧��Z��bO9>�Z�m\D^%���L.�y�h�;����bv:Ѿ���eJg�n�����j.�3�Hu,���>?B���B�Q)��\
�WD�	��9�D��^ �2"b��x���� Q�&>{sLx�M	*;��9;:���ҙ	��t7ή�ɸ%��Lޕ�����P7U,)���ʱQL�~�6���B�L����ߩ#�)���	�"�kr��R�*e{u���uh毋im��r��/�ZUӨp�	t��@�ow�zlG���q�;�\��℉t��$ ������E�piFo-d,՚���7V�����k���8��|���;���;/}o�$:�lC/�G�w`�M�I����K�U��i��p��R�q��8���-NQq�j�@���:Ӛ��k�P������[��c�Լ��An��O"pR����p����i�j��8I�H+0C~�R"����Lv�(��';���E}42�8	~��kb6Ģ���~*ш:Μ��gR�LG��u��6Ri�C�L�zJ�|��Y�p0����(�A���/2� �I]�c.�,Tf���2�{���}�8��a�,TZ�����x{9��uqB�)i���ӊ=cD6�{�Ӂ! ��J��`1Ȭ�'�k��EN黬�U��DL�ٯZ��Ѽ�𩗕��Y@��7�U�&h��w� ������Y��\F�,	0S6U	S6��$�2e��N���"0D).�fC��l��y�@~Rv	�=�q�7Ů���N�}Y�����f���A �!��v�y"�
�n��hXqa�e�n�~��u�9_O'�I��$P�XV�]^`��ހ��!�"?"���7��dET<��άD)'u�_տ�Jy��{���� T1�oo�l��&0�O�ǐU��J�]�!����q��?(Gl�:�7D;<E�x҉����ډ���t�۽I��N��Iaٯ�1�uĲ�g�D��ZRF���:q�P�D=.�$(�ܳQM DS���U>Bϥ�p��M(A�߉i�r�^��gB��르���� ==���B�۱ Y�K)1jzP�ǩQX�Ө���V�����%��x6���zx��v<�#��H9;����ݦǿx����Xԁ͖���&�<@o���@�i��D_�H���
�'Z`�xK���J �}����Q��	�Y��I������%Ӄ�e�U�a�e4�9X��"��R��>������~.��3�k줽tqm�c�������v�&�ۜ��6���j�ZG�Q��g�B)�"��<l�RG�����HV�8 �̦!%�})n,q�H6 �D�����N��R�_m.�E?3����8q�?�\p*�A��&k��'��W�%:��r���(Y�Tj��%�[���1S��v�S9<�F���������%�w��c��T�(k�nU���J�)Tjɛ�6�ʽK��8�L��IjJ��#L�����c��|k�"Ů���1D�В�>�Z���^���� �6صx|3Ǥ߷��gc�^�f��١и%��_�ͯe8C�pw���mF{���+
A��^��}O��&1%0#9ڦ��lF�m �h�g2Kxq���a��KdQ����_h��P��Wio@��
�Ws仕��_h�	�Q�#��Ǎ���N���j>Bl���Î�	\+�rQ��tTf�)���KG���]!P���)<a t{�R�4#�ZSj��%K�OU�7rIId����<`PO�L3�u�"�s�3RlOI��*�zxsU�Xd�e��|!Q�7����7Ϻ{��^��1*��O����[La�-|.�D�Av���خz�X�6v|�o�,�76EV�TW��ѕ�6L�h��:�b��s��	;f6��zV�5�P��58�T�`��_y�HL�$TA�tUm���"����7��!�����M���x��m��Q�D�L�I45��ݧ��W<Q�2`����g�h"x^�A�j�rfJw7�(�J�IOJ������o�x!<�R�3{{e���]|!���-b�ɭ��U_�8{��d�ًM��.H����E���:=T?y,���j�����H� �wC�g� ��>�ɞq%�ە���F�g��uuG�gM�Q�L3�O�)�$`�G���o���r�c�dp8�P�|�gF0`n�=q��&�9��G� N�3�4!A@�|Y��^��/�%m�(Ӯs�Fs[�)T�"L<\΋���hy��!����(%�Z��[� J���"�@KVK�Q%!�S������x�&�s���.R����Ц�mo���p���r��Q�K���<mh �Q���?���-�*���G��Mx����C�	=0��)iy*p�P�k7��ηt&A�9G�m~e˯Z����&b2q�(�"���ҎܪkZ�oy��\7(�1�BJ�E��3�ckX4�a�5�^N045��������\�y<G$�#�(�˲ϙ������1�P�T��e�� ��K$�k��kH�#�ߌA�m�e�i�A��&& )�Q9�L�N������C�-� ����7��|삗C��b��=2�0o�����SL-G"���_�M�h+脆J��`t�WX����x���&: T�i
<[c�I�_(l&Nm�uQ��!�/�!�}�-f�ч ����1�b�����by�xF�"�
k{�![$V���D�8^��/���pK�3�#���:
��ֈ�"W����Qh"���G�x�j��:]�t���"��`8X�:�qݫ��#`�"}:)-@և��v��>Q,\� k9Xx`�݉ᰊ�%��4�w\pla�U�S�g2G܁��ݠ�|U���󩜃G�N[��v�#+ߣ�0�/"'�Es)?��H�z�G�1Ia���ߓ��K�+* ��̖���5g6�˰μb<�8a5��^�2�xy#��(Q&�{Kc�	?i@�����4��6��L�p�˲:��d��wD  �٥
�Lq��gH�P\���Vݰ�L�Yeσ��<*�憻�G�.�P|	E�BΫYf�]e�H�T@�����3�k�����v]�E#�����j���Q�$@��\��F�:'c�Sp�*u�7�]��,�p�v!8a�J�`�y膟�=#tl��P��w���,�/ȣ�������~�ٓ�����[C���N��/�=?�X+��wQ��:_����,Vo#��Z�u�y�D	P^2|Bz��dw�����[�b�1<`ڿ�-�J�UҢ[�m?�w9C0m�[IF4K��'��o	I�6�*>� ��'pE�ݺO��Js�K{t�	��d/h0�
$D�ǂIj�N�/��1�_�w��?cж��u�U8߹���k�A�Q0ɱ�%�K�'�pҴ�v��JJ��J0��s��J��W/o="�[e�WQ�ڏ� �ւ����m�i����#O�<l�Qv�y9�����A�Z���S��y�t�����I��[r�G
	��X~;%���&�ו�]���W'�-ɒ�N�z�R�e�����`��
Q������ސ_�F͚�J��T��)�
w�jf��uE\�[��Q8TBZ(��-��{Y��Ϋ�Z4�1#�a,�����1Pׅ��=��) 5Ĩ;�0�v�w�މ�޾�Ǽ�-��n�'�ۇB���I����>-� 3�# �wg�ʀfBLQ2�dfՐJ'�$T�+͡E$���(�Nve{�O��`�ǡ�L��8�[�/F���k�=[yjԶ� T�������c��ɕj�䔜C>�k�.}�����i��j�_�D���M���P�LnW�I�Ȋ�H�l�PH�H�[�f�%ꂽ�͘N��>��]��աd{�-2&�5�#v�`�J�4�|�Ѻ�U�����bt�N[�	Y��x�z:#/��W���\��ō���;+=��p_�/�,[J�����NҨ$�������p7���r_��A���@�����ƨn<��2�z =c�z귏W�<��b4����M~ήeI3��)��N9��$&�s���{W���t~�
Ԝ��-��)1!Śc��a�b�|
V�>���5��߳I�%�y�
]����E�@CU5���`rF|�@f��)����Lh h/�$>�|�D�`_�jv�L���I4��Ե��W�C-�lMB�_Tq>gD�p64��P��I���f0�ޤ�L�"�f+
�ȵ��_O�G�0�'�*Mtcv;�~E}5��y�Pc�k4��hP;�V�����,�[օwƪ�5��!�s)�v6CK~�?I9L���cޤ���H����1�"�e�G����k����S4ᤰ��-A�����l�#0��T��]�9��"��}"�X"��-}n��N��X89�rW���;�E��8�6�s�9"7d��z��W��}� �B8_�Ȅ�uo@O�O�� w�5:�<`X�B!��_l|fh�7��P�#%�늶9�tؒfJ4���p�|��;�U�� �����OEl�����ȇ�`3��-GA��z�@ 		��Yi�%��>ׯV��9�����<
.g�_lK�����p����B������j��>��X��K�E� R:���G�㊂d�����t^���ퟲ'�</��`�x���Ù���|�g�������P����h�ֺI�q߭�+��i��y$���Hb��ky����S�*������2c��Acq�G�"d���w�B,ϗ���q���TI/f����\��i���H����{��`�X0��Fv�HN3�Ϡ�񜞨{y��_8H:�G���o���i><`-v�S�2��ъ�|��;A������ګ�����/�.s촐Ĕ>w����!���,��|�Q
%nh��z��r������p�x��x�>����6@]����[BH����A�������}i�@�Ȩ��m<V2�csw:2;qj+���:�/-���݃D��?n�:�Vd�]�|�?�,Ʈ�)q�G0HIL�Y��r�o_s*�%�_�[b�"~K�D��Ҟ��`|��e�<He�')ttc2����Ξ�gbW�x�6�:��2�Sߎԑ�����r��s��!��H
D�W&�Ejf�����ڹ*	�h��z�0ښ,mdTADѝ��Ֆ4}Ξ����,ZccpW�8r��'ws����W{������D�VM`�[�yx�x�Sx`�P���]�Ȣ#f��ϖVɊ�Z5�noL�QCHũS�.��|�1���y�БTm��n;�����l�9j(U�\�$Y��>hy7i�5a1dP�#��-�L?:���a$��Z�����ߞ&i�'�;<Z��gF�3����#���20ɂ��KRi�9�UCc�=���a�+�������n�;M�Z��N�O"��ܙW.8\L�Gj�
�h�lǅ`��1���o��;�΀Z�f-�Hs����U��um��e��"�71�I>pdF��tQ{Ar![����Jx����p(	0Í���w'������e�����?=>��J	½G�_��ɧ����g����]<�{��~�6(�{ZnD��mv��<Y3�����:��{$��xz��g�YEWB�I�u�);i�}�1�E�0�;�J�g����܀"zB�^N�mm=��)�l�J��;�,.7����U)ג�ч��q��ָA�C~)wW%B��+{A���l�u+i�����b������-��Qե����!��_��-�2v$��5���l�Bm�e��z�|�97t�B�c�/@=��n&�����������!�Ӛrj+7Z�P�x!����S;2�T����m��N���%�7	� .�D'��*:b/�`���Ȗ�ǘ�4�d���3�9b><ԉ�ku���!_�cJ�#XШI�E���;�K��+� ���Ux��!���2LE���ש��}�8;l;��ow��q��ڙ���bB{��&�.��هU���ټ}��_}��h�-�%1�)�ë-��ɩJ�HBp/�g��̥m�͐�Ŝ�28n�>ս�U]�#g(��@�J��E�z�� �������A�a�X1;�5n�=��T˅�U�D=����d�L��p��B`��.�h��i����M�^yHRQܲ!gc�x]�`ڝ�M1w��/�x0�+{��gb�Խ̮,�t��X�?>t¢ޒ{�bې]p����k:��C��ƞ���]ogU#<f�xK�1j�ـ���&�{�Q����'�;K�O�3>+s�����=i�"b~&�M0��a�u�fw����!\#p"��%�5u��3�$�-�|�Q|���0��C���0b&y!HP���zB��{�P#�4~�+�{�i�A�9�������2�T�҂�5�-��:H�it������'�w&�m��ȫd�����&/�,��JK{�*��n7�nW銭Ͻlmg���$�V?(����V��e�o����}�I1kXi�Lҩ=fo!t{�l�c��Tq,�e��u-��0#�G:K=54���Y)d�lW����<X� xC?(�,ކ��y�F'����B�M�,f�r4�����7�'���sg�	�O킡`eh�óbsxQbJ��m*��㗖��f��7�m6W�H��YI��D�>"-�퇵F�B�r�Ҵ�F�f�L.(#O�:�!�Ģ�1�V�f����`�E�2hT��o������dR��0�����^=�Ҽ��ŲSte��h�����������ٌ���Gu�2��#��) Ev���Ui� o�d^O����m�5��CY��O���\��6�B_>��Lߑs�9�'F�X����+��G���� h�X�����Dg¾(�{'��X�A�n�ݶ����|4V�NG�ܢ����4_�o�R��ńk�w�h���RҼb�J�ɟ�:���tyw2;�	G1w���Ġ����X4c��y��l�5��5MA^L[��o����;���	ry$u�t�&�_�d�h�khD����-塗X��]^�I�ȓ~Pa��Ū�d�G���\铴mc��_!q��d��'���m�AK�|"1q����$��p��տ
�Ir���?�S��uj�*9.��0�l"-4�
�Yg)8|��(
�Aq޸���	���7_I�X�v|��O��s��!���I�z��f��#N�,�$�DP������@-Z��Q��)c������qp��$#�Ӽ�
�D; -�e�Q	/����������;��H��!��J��Ty�(�0����W���K>o�w4��y�l���d�/�~��x�,�KݑP� ��]u��KX,;v�Z��w�t浽�����y��]?w�!�7B���;I�w���6 �ÑU����[A�i�#��� |6�!�n�%��wG!����%�j;P���QzQޒ�t�?q[����8��Z��@���X����iU֖�7<��J�
�����%Es��Fq��0ܰwG5@��܁3�ӗ��b�L�&*a��.�LT�5�
����6�ԉ�n��/�v�q?!>�5c��C�``a��z��뻟���O3Xߢ��t�T����ҝ�jq���&P�c*G��_�����P�n�o�KVn!֘aZ��X���U�I�@n5���L�G$���&���ɛ�m�z<��bP�vBvQ��q9ldW����p`y��yc}�-�+�
=
H{9�<kmQ눴B�Hwi�)!?7��E��Ԩ�oK �&�=�'��k���y�~���N��v�!Aն"�F���؟H(Կ��/Ek�>�z��ǯͨ(���ߛ���O�eV����:
�n���#>�?����4��!�vW�}�c�W�_*IV�^
1� w�	2�ziD�W��Y`6?�Ῑɍ��y�#������?�:=S]�N��4�����R�r���y;\��8w?䩃1���rx�!���� ,uܜ��!X4��;f�\�F��� I�s G$ |=���_�ф�>�S�:d�+Z�$Ϊ��6Z%@�8'��-�I-_��X��W7��"6�fz�ɼ���`�QT�?i:SZ�������g�7�3o]F$'���e���}��fX���đ�t�O�z��I���,cRd෨!�P��Z�t�q�T�<��N��< _�Ë�L*r��a�Y�� u�|q�\n��z���|'�����X�&Ĩ�{���yj��ߌ�~����f	`L]���)6|7g��}�W��o*n�������M�ÛsJLђ��pR>�f�w6v�m��)�8���J�#��0HL)�HX�cQO&�}1��,���k _z�4�v��
^q������?��sz�6�I���♑iEoK���h�W���qLڜQ��NתE<�_kQ2���=&�⛆Ps(�l�F�3»�!þ������g�a��Z�С��h���
��A�����n/zM�^*�z���5Z0�f2���x��Q&��bT��jfG6�]�<�F��bs渆}DЅ���y�f.ɔ�����F?Fbz��-���5��2B�T���t��t�_���W�0��n�QA�j1h�s��E�G��׹�*mÎ�����~��:O�c�\*0yH��v�',��d����k�LRr�7��~U���j�?��e�'t%`^VM?�ilx	% ��D�I����1+���6��=}$κ58 hz�}�3�;�2�ӡ��N�7t4;�`�:x7�
���9��I����+lo-$�)�~����K_�`f ��G	���2���e�S�1~��2�=�ͳ��)��hm�;5�S}7���j�K���%�/~�଀v��+ѭ�I�/!Z���+��.�J�D�(�ĂV\�4��ރ�����#'sKd�����;��N{��7'$���o�Y9@L�EW�7�$�{��ի��e�%��q�e�@B}�%�����% ��@�����:0�8U�E�x���ꭥ��;�z��M�3���BK�	W�G���d1R� ����a�
�v���M0��	����g��N �sQpO�����d��ec�%�;��{�<�3ﶮ,�r>;�q�0�͖s��b�A;�'g!��3�.�`� ��T���XX�:y������3=�|��	k�۷xN�D	��91�*�p�GH��7ɀ�!�!g�,2mr��<�|Ϸ5�,�D��ar[x�ǅej�(�guoz����a�����;��r���!x�����$�h�]vy��Vc<2QB������K3����'ֻ�c�{��s�ܡhc�c4���~FS|��O��5��O��n�7]�s��+�gR�4���)�������X���&���{�NE0���xG��*�I��u���:�q�B���v~Qq�Vm>0�+͡�y�i56��n1�����}<����b�����9Y�t-����tA�z��EF�M��t���9���7�H����}<l4U.,K���G��G�{oܼ {������@Rr����4\�
H8�Y��x�ci|��O|���8OS�p_h!hd� !ܖ�к��)۫��\%<��S�% ��X���~��S�Z7�~�5�a_��1	�M1\U.�MK[����?�����J��X�~J�!�p���F3¨�]]! �Qʏ�☢��l������hNR���-�=F�qN�w�Uu��I��]����P�1}�����O�����R\����3�wF�8�k�[�[�@�R�\R�#e���'|�l'����@��n0�ʂ
$d�fw�[�5���ycb�#�& y�
 ��������yG'_p~�24N��O���2g��\�L�Zq&$����aݰ���{�5U6�;�Z��8��� ����䷇��\�b�\i��ԭ�G_�b�~��-:�ˋ�� 
���Ԣ%Wn�FF��ۡ�nqe&�[��t���d�D�J5h�h|i�����,3*�����.��3�7h>��������)��0c}�w��
��u_��A-߼">��^~\�Wʚ��(�$�e�ߚ#�f�*���d�W���78��8�*�IU6Q��Gӆ1��������̋�}o�%��}_��A~�N⃂1��*++n��ȦU�ʭ�k�`��K�
��9e���*��jp������6������䑲s�0v��A\%
����+1��?�zmcH�:*ŵ�k�h���f&�Vl'���
�:�1[{+h��'�!0�|<w�W�Jִ��wZ��{�3�h0�����7RN�Za��ab>�6�M@K���~jU����ʗ��G��	��3�qj�P��.�T'��Mնi	�u�·�o�����'Q�@�yf/�f�k��y���}q��#�%u�'��{���zH��={�*X�n�7S�{@=2���޵U�(O/�L?3�!;>� �}�L�.����y���?O�v�綱��:]<\��g��#T&�2��>�7s|�ߏ2�f�"�~���(��k�l�~+�{Ó��5e�����9�ғ���̶V�
yV�X��bUMBU���.���8	��U�U3 �"^nu&/�?�
I�u�����
e�T|�5���+�I�Vqm�(�زZ CEjC�5�Ј�-|�T��h5���~Ro?>U�T;;&�z��A� <�����M*V%�����* 7cY?� hԠ�j� �]��֧^��Dgp{>C��̼�V�R�jgy��]ˊΊg�2�Aآ�)�TǕ��X�a�N�A7��l�?��%�t� �2F�^C�Nv~x�����`�1��C����	;a�����0�>q��]�	�5�|�-g�Ť]� 2?���ˤ^m���W^.6����X�F���%�Vy]m-�N��SKӻ��*�4����9{��B�L��Vy����T�3�>\(�z��+؀�E��>sxu�e�D����ӂUK��L�Z�2�Dv-�l�d,~Y2����L�+���K���C_�瓂��FR���"��te�d����̿r��"��Ic2�F��Ʉ'��C�p�u��);�$��>i>�X�r�Uc��� _�5<�By,w >�M���T#O�F�����A-Yk� }������+Ի�@1��d�L��� �b66/N���H�Ђc�\:��Htmκ���؏���T�ީ1��#��<�����nm|ÕI������FbY�]�Qn��\����ؘ�%=]\$<�5���K����
�d�R\�hW7ST��i��m���y;�nkA�Q ~|%��ϑ;'d�n���W�����Nd�����6�nOu���+�'>px�A��5ڙ�.���\�>��A����{WڧR�`a͏"�i�RL�N(�|e
:�Io��j��u��AJ[�l��#��D�����;��q�+Z�ګ�9����2S��j����G�6@8�Y�K�ĳ��2Nb޴�T5:<T[�2�U�P+�Wg�)sX����'�� ��H����#N�����1�K�,�qL[�$����j.Xl OwO;5�|���]^�D�d�֛���$���喿�[hV�e"��zfA:�׃�P���ۄF,m�kH�&w���bZ�X�RM�Ø�EoH�=��t�uTI's��K����Ȝ�I�`O�#�0�4	��ɧC���T�ty���FΠ,�B�]���Q7�'AzhU��~�Uάɴ���!��o_rd]dg�L��'�lOAP(}�7?a#�
3"c78t~a[v����Łn���^T�5J�����uhb�#��72�>*&5.��ضl6k�')uzO�v�3�"�c�X=��u�!��+�ɧ�sȕ�p2eޏ�滔4��`�& ڲZ�%X���}�|��\�;z�,��̛ܥ�����v�s۩5�{I�n���No?�!���/�UQi�������'��X�E����v��}%�(�}x�˔Z��h��l�ϻ�R\*!s�3f���<��mGb�8y$)j�H-/�^��<��s�XcjH����c��
�K5�
_��O&�dވI�۶�+��scyzy��D+����L[��t��"Ҳw�M~��4��Fs-4��e���K�:�S�xTԴD\�z��	ܗ N���$�ٓ麜�XL���2�n��_�8��C����.���\�(�U閪�56�
*��+�%l���RP;l�ބX�b�ۮǴ��+�_����Z��#�!u�s��\���c�q�Yf-Բ��T�躩0p؛�ks %���'}9�1a�e���M^J�TK&%:�P{���d�"�����.-,lB�jN�	��I��^h�V���{?t"�n.b�O3n�����n��F���$�o���Ds,y)�5�f��*��~QimR��?��#�h��O�⾥����v�;Y�R^��GƱ�fcJ�@1��Z���u�gHm��f��}�����d��|qݓ�ؼl񸓌��H��l�pkT�FP�Ə��="�-�K�c�%o))�0ڣ::����e�������߶6ɥ��0Y�E�_�&��/�i��A%i���\'3=7��n��-��C$ؼ�DK�!�?�x����{�G�SȲ�G�����|/u/���Ք-S1�4���ي<�\d)q�U3�ڹ��"t�P�/4}ɏw���6�}� �vƟ$�Ę��=��ꑏ��)x��N/�%>I���x�IS���ӕ���
�����̳�4,��b@�_���,s-�lI�,x��uG�R��QC�uS����5������bF1m�����9 SO�ja����;�Nѡ����lB�x��2�N� c�^��ׁ7��'^��1"��(��H	�m��i��høJ�ŢZ��cZ<)��X�II�_����a�M/&CK���\������������I�F(�f*f(��������BTmO��?^��=n6��}�p�T.���Tq�[7OCD#(.WD(�"]F�H��K��ӣ�{�ny�j��$���=h�֑�p�H��?�K�"�1��
�!_[J��Eq�,ۿ������V����~d�q-���J��@_�oiT���w�[�Ƨա@.$��@���m`�2�}��_�q�^m�	u♤Dl��?��ā`=�sZV&�ؤ�hdSq�X� 1P��%���3G3� �xw��$�4ft���G!�wE��-�y>Sx<����w\��t������H�y�wg��Ѩ�mCY��Bu���K&�L�䳩�}��"�"2]B7�M8/5
��Nd��nC��H��0*��]@��R/s��$0�E�H���[f�9C9)b=���ۏ�H��X�7jG��9�N�J�.7��}�&��/D��|4^����Q����O��&�� ""0�kƭ���
�[���' @�^���]D�bk\j�+E���*�\ڵ� ���;xA*��"��� AI��Sv������m��j���:�7J��{IA��G6ߠK�r~�����=�_�]ĭ�B�|z.�Kh���S���!\E��� ��|DL��v<;��1���cM\��a�EvG}�0+�&i9n���S"���
�Ie�f���G/Y�ib|����:�:�g���mYv`��4� ��'����I�ۘ)f�ؙpT�Aլ/���#{L΀Ak�ݒr�<�灥~d�|�eT)�h8�v@K�'M��d}|��_��n���m��ˠh�"��;~ʯ�>'E{�o�kF�9�	���2��H\�F-h�?�$S��J�-I�u.Q�]��jbKR��	`�+z� �鸭+�]ǫR4 (�.��R�+����k��
��$�������)qr��E��X�����+G��_c�O]�E���*W�E�7�	ӡ�a��@.6������ x&O�F���P��.���W������'U#�������k(g�~�Q��^��+(�ڊ��Z�<HRT5�r*KɁg]N�D��SR�����`��e�ñ�k���Se�&�L���f�&/X�Qa��\�
�r�
G�%�WJ���~AMl/��� hFw�G������� �2H�ÅR}��h4���]LiW�s�)��'1�F
��R�Ǝm�㢴���ĩ��'�{�h2;^��w���2����SW��l%���g�X�kl�x-�{�+$�3�U��o>�3��"
ʽ�eYG�s��IG���^��y��u��9" M<��"L�5MJu`��(My��:x������m���d�ɉZI�rZ^��{��R��<=���	��/'=��#"E~+�e�X0�sH}c`�n�u���j��Wy�אa�Ό�:�_�*~����ZP�z�%<dᤄG��P���db�q����_bI�m�eAP�1#�{�J(�`b�1�bրo5�fb�3�Ǧ�1_����7��jԞY]D3ϭ|����L����R8�6��m����	q�E�r��(�W���K�QD�`������UlG*s��v�nHܛ�%�����ؠyM�Ɏ?OD�Ö�y�[;�����|��'6g���Ed���mnDT��щH^d�!BS���QK0 ���Xl6>a]���a� r��p�V�<r�A}G�|��~����.0�2��M 쫹���7"�ڍR���u@�6[a@��nھf5���~x��E�u��}/�M�&s+�w*7��ts����~d� � �q�=f��Ȓj�*�a;�����ۥ�%y~m���y�ކ��N��yF%$��N��!;?;��X�'�a3��Ӹ�?9�2M��7L&��iu<��ǒ�� n*F����"�A�f�%�\t��M.{�9t�M��#�^u��]����l���ꋫ�ɼ2T�
�����G)�/:���A`�����B��)���6�e*ԉy��C� �~\Ҵ[�Ӫ�e�{ʟ�%P�N�'(�k��U��;��;P>*$�?حE\�#�&�R�-�_nɺ |��f�kKY`p�q����irs��l�ӑ�c�A/��E[�D��	}��e�P�	P\��UԴ�'�K��TL7'*�pj��2��X?�����3m�,�[H�������U�33<�L؃ŀR��ѽ,�綎�W)���`1O��/�W�H�Lx��,�cX��$��ޡ����T������*݆��CF�_�pbE�`��V�SUX�J�q�qyA�CqsF�If���9�����.���G��O����I�RG�&�O�v��������o�m��fkA s���D�{�L��Yho <��	d<]�^��ގ�!61/(�M��!���ʿM�?�3Z^j˫�:�3�^���Zηx�ʹ&Ui��bsA@��C��,�.$D��?G��[���&k-�S֧�|Z���I�F���s�6`3�}c3�eW��E#�~`��@���j���ii��>���8�DU���M:��f�rzR�Z�w�����؁�b��ؗ�����5�	t�ɔ�����Ş�E��&�/��@2�(�3C�i�~7�������t.cm�'� ��ɏ}�۽�[	����x������ܑ���֒(#0|�B���necx*<���:����h�=����!=T��j�&�D��bd[YkY <R�Hͳ����4�L��j���}J4�e��n�#��"zͫ7� Rd����L�H���M���Y0S{Ӷd��@<���}}H�hH(L�cĲ�)��)�	�~����U����F�����\��Q;����"���lT���-5��ߟ�s�h�A��r���/�}_%���b�q����'�J)$��- I�^B���\C�-�'�$�)E�+~#��g-Fؖ�i��?Z$(z)!�X�l!�ASR���t��VL�~v0x��{���-�G6�u�#c<FA���j�V�$�Ͳ������6�� s�ca��~���(4Ϊ���w�}��P���yT������ ^���J���%&`�"A0���T}�$*�����Լ���/�]�{ɛ��5���o�~��-����\du�ʍ�E�}�y��-u������R~p~�'�4�/���z�4-�F�� |߿�LE��d�ٲ�%�"��if�#gZ<]J�aHWn�ST�%�Q�+k��hj�9��`�@}�h�o����ܼ����FG4!h�rsOZ����6�a�g��)m�)+1�AL����6h��	���#������ h�0�0��Q���US���wv��'VBK�p�{�ʏg��pl&�d�@��N���k L�lj�f���῱�<�Y8�<�d�@˟��u������ߖ�s����*m��(��4���&�u݇<0���M6~�+�#�I[�3��ق�!$���[��v�V.Ʈ���f+a�Śc5]1����>�I�4���r/���ק��iYhlW�����s)a,�S��/�@�y��d7�$�xN6@��xh�	�!$0Sd�@���e�#`��3s�l5%���:]��8m����S�
u��1�\B�PD��'�d�,�������4?�{1��R�'�=�8e4��Q�,��������\�c�!.���r�Ď��=��nr"PO� �m��y۪U%5�g�E`��ݷ����V���^�v��1����nXF�=;�ާ:Xc3>�4�,et_�m�zD�T�uGV����eF�.&�L3v\��mڠ5L̙)@�K�'���!���Z��;)MF�����_�����aʂ F^?����=+�z�3���>�ѝ�����Mn�\[U�.�l}�a�Ҝ�-4��������ge,���-	��91�����,�UV1M-�`�]��ƓG��_Zb���Z��?�hd�;b�^�:�N���W�Q�3�Ge*���}�r���9�,��˚
$�$����;�Ȭ�_u ڮk�\���y��+~T� i9)��s�iFl�X�x΁��R�G<��3��ez��l�B°R⃼ ɐ�<7���*���E�a~�u�2���T׶����d&��/5!��w<����#�r���r�%��i��͔��s*9 O��4%;���*]��*���|u�!�\�.
�݋?�arٶ=�󋛝����9u���gќ�'�m���s}�8�������p�d�����Rw���2EhT�6�ayb��a��o,г���������Zx ��|}MQ����;:xI�|�.>2e��x\бN9}����,<�4Dx�DՈR
Z�X6��C�*�C�l���>���������	m��%'dw�Ūn�g�LS�:�a���VJ��y
��%��w�T�U�0|r��}�OA�Ij���{�5f �o`�ו2�A�?��7n D|e>Ĥ+���*'�븡�r�Z��aOg�w^��jn�,+1��>�km�eQ����	�ٲuE�R��U�B�b�Y�J��1�Bqw�e���+1��S����o�����_~�$��]�� ����Nq�����8~�<)I$���\�+Aj����[r�+���i� o������,�̈́��o��:��c���S7ZZ�C��C��m��5�C��*��z3fKNK(�{�/�m�1K�FIE��o�i5�&QV?`�e��kꁱ%;���ا����?����:��!�:�#�ߠ��q[ϔ{���s��P"�u̕���"2'4����QZq3P�$H�d|# *Ϻ��G��%L����cA���⪳�؏[q^�m)D�o��:ME�Y�e���M#E�6��[�'bU�Hܱ��n�\��?2�E;�:�'9h� S��S��7�0V:w�6NҰ���:��P�x���qaA�ZDz�6?Db۪MXiWH���J0�պ��Y��Y���姮�L�m�`\Y��7yP��j�Dʹ`�ӕ�F֒��q���;sz�N�5�mO=A2e���Tv��x6;sj��|3���=�����C����큂HL)��B����P������)E1_
��F���K$A��t���'L-[���2�~��,����Ц~"̽��ۓ �?b�bBIߚh��E�:}g����Ē�=ҿ��Ug�����#���鷵�nR���a�*����h��&��ЃWIʌ���9#ɠ�xL$�yħ����$�L�x��l��p�^��d_Tٻ3���j`��d�o�'��3<i+M2�H����(�{-�A��g]B�3��mn�e�U�H����7JM��Ɖ�/��8����a`kXfր��BD�0*8v��:��$<Ղ~dV�OW\���Ei��4�K;}%|
��^�'5 x@^W�gb�4L��O_|��@���0��"܆��7�R�:�cp�p��M�F�UIP��s��W����FX����L���}��W��/I���͟���Y1--�\n�#��g䷯ڜ�B.0L܈c�Blzwc�;��x*�(�Av�9��*|: ����eԯXPz�ܱ�bQo�Q��!���*>5�O�o�k���:�i��$H�@L��D����z�hv@�%�AQ�I�����z$����੊lͩߖs�4>E��� �Kc�!����Hj�Ь슲0Iik�:�o��S�L3d�RM<���ϟ$3��&n�/Ss��/Y�D���im&EY�
v����ö�5z%�nص����I�J�ܔ���d^yhs�9�,m��<��m1B�<��9���[g�(.����Xҿ)-�B�{\�|˶F�t[� u�����+�}'a��]��O���A#�����!��h�:dٸ x[룰�6>�8����u��T�~N�T	U��_�q!D&쓕CQX���.�̠�5�gmw(�%�W};�h�	֐�	�9N�M�k��^5��K�}�Ό� �"����5�F��Z�^`YNE~F�5����8'�x�$��G��1yq��f��_�+���L} ��X�Ld���;�׾ܵ����s.�� �����jx��6�6�w�i)�����n��%�[ch3:	��[�x��Y{��B���*�Ci�	�������\��KN��r#�!��^v���)�p_YS��'�S���16�3�P@U�R���6c��r{wE��]]1�Qi��78�"@���!��������D�i}��s��k�������}��q�%�D�Q]HDL���s�n��t��N_7]�j�L�@$G!5�d�@] �����+�L��)� Ĳnh�h��,�$��%�1�?|^|�E�=���x5��0P�<���R���D1��]+a/��E�gm�k�)����G�+�˫5�K�H=�~�,)#І2.��X>�z����,p���gOt��9��D$ݖ��Ԙ�@ζ�yy��l��Կ�:p_���ڛ��а�_�D�ef��x�}����[b�4����'\���������۸�H�e!/7
Fbs-�;�_�A��r
��=|�Z6z���3���oL�I�F�2%xG �]}�@��Z�EH�E5Tz��R�Q�:}~�����X�!ET$щZ��|"�w*��8��f��b��j�L�"�M�3!8B�C�{D�3�� ���=(1��x@�	��]�OlP�0������s�P�=��ù/�E�a�^QY`	��Ⱥ��	d\��.h�����7�ś��������;4�y��ƊB���W{�1`��Qq��d"Kjr����i����c���,2�Q%��p.�Zg�e�t�m.���^Ǵ�f�g�v[�M��~�)�
\\x���Z��*N���[Ќ������^�;�ݢ�m0�prDe��2�j\ex?�f�:����C���K2���ҷ3/�
"�q�
����&��ZTH������"���*��&�{��w.^~�m�N}~�����_�/��[��2;��fI�Ÿ�W��Q��	�d�`㰺�� _##�P�hぢ7�pC��u1�;�0FƱ� �؟R�Bb�,;���~�fd�S�)6�@��A�3�e���f�3�y+ik�0�]���~�~�@g(B8D6��g�h����)�OH��e�e�8p�<�Ơ�gѨ�ɮ6/��Y0lʝ��* ��9]�3~�A����R�#��	aL��@U?r[��M�4�&	o_�.�Hyet�&�o*����5����EF|���q?�4,�L��v�R^Mcw���	�h|���E�;}`�=ռEƇ2F�Ru��Y� 6�z78�Xƒngȿ?%�p<A�;�%-(��������+��>��NV�F7Hs~FJv:􆒳\�LIT/ޠdjx��91'f l�w��|>���o��5
	Mb�� -GI���d+�a��F!�<D!C��Jc���2Q-Bt��䚌q��5�,�m�x��/�K\��a�̢��y.e��筱��%g8�3b]���S���c �	��~lo�B�w�|� �%�گU�!�[��9�|J04�l�X{�2G!�>˟q�\���j2��,fx�=X�-W|ָYPh�\b�`��Hr̾�H���>��_�����O`����{���.��݆}~�r�7+�!x�ݦ�>�m�{�s<S:����)�������^��) ��g"�~�:{ o�Mj�7+C���,Ġ�/F��S�U��	�J�>]Q��7E��SJݚc�۝oOCe��1�6*fc޾���ǜ֤�Sh.r���cq`XY4�D��3r�`���i��������!��Xa4�R�W�'��V�α���JܴNg��a�cw�����u���[�X�>(�7��"v����dim���e�}��U,I='������9��huR���D����M1p��Z�b� �3_O�l<`Ν?Zv!Һ��z��K�(�g�����e��R�j�[�*JM�Q;�\�,�.WϏV�Zt-��
/I���Y С�#`��j[%���6�se�^��h�ܨ��`�f�U��3������K[��XƟH�Ţ 5'
�a�XW�du�ئK�QO���e�>(�o\@�l��/.t�̣ߙ}0�
����ѵ�[�h(�-��L���#�����A%QH+��ٺaLU�t��/3)s�"x��j�w��#�FN)v���*s�4U������5Cv��G����E����DPA�c�*PC��`~s[&L�:FpN8q��Z������PSC�Vb�6�B��4�>�z��n����@B|���5O��D�&*�=m�z���9�#��G���L�M=%` Y�|����#����9xrQ$R�-�]؜��C�nC��E(o�T�
�P�8k:���m�B��g
]���"�ܔ�7�y�����d����	��`2�v���h��$K�~�G)>Sʺ��g�*׋+#��f�V�䲠ӗ�IЭ'�phZ2�Պ\�1�񹰟�^����2��������Q0d�㺓��,��|~пz�	n��[!��������F�	������.L��Ǩ��Q#4h���$�� 1�J<6H�'q�c��iZ���'��q_���m�/u5v�΋t����J{U��&�ឱA�𐑞�,t�Wm�l��v�lS%cGãS�~�g6�0����,�RJ��x���J�x���2 �a�KVH[^Ö����lq{��b�
F�f�{�d��'�I-�j������!�CqR�'���<4��F�7:f��*�]?��+����|�F�4c�n��"�u3R=�1b߀52�"o84��J}����*X-����>Ȫ�i�����p4[l{ ���
����9Va���f�V��z��bv`6�9@i�5���&��p������Υޞ�k�2c�deoF��������{n�^_�u�^%��/I����W�Ǫ̊N����n<0��?窅y�8ZC���mi �kr��Y�W_]�PC�c�j������V��MBq�S~��U�ߑ��+��%<�ts�2%��*�x�)B���|��bфۧ��_W�v��`�amE��<(�&Svz1��?/��	f3��}a������ ��d)�C��	ݜ���U��̙�~�g[�jM*�9������e!��:a���L�q�/g��Ջg���=1�Y\�����*�A�oO]߲xFDrQ��+������{�|������<'t۳�+u��b�������m\6�(�2�dM����M&Q� �!�����]���2Ah�90����~��B;��]I�2XSE!���'t�]��(��\GfE��zi�΄�prM���=1���'�U�jlm�i�&u��sLՋ�j�|��I��0âW�bJ*� m����QI��������}F�	��(���	{�����ܦ�Q g��� �'���/�U�
�ɛ��nك�g��)44��M	����C�`�Ya8'�켺� �Os�v�}
�L̪(�6*�(��΂w�)F��sU�HU�h�����}��UE����2���a=�p��I����m�-�D�{J�ER4,;���3��xav����L���g��4Z_�E�R�ӭ�rx�;���.ۊ|�����2+��bvࠕ�5O���ٶ�e��[��z�!Yj��
�I6�]�Pd��]uS�,G(�m�s7FrK4u���/�i��/t}�~�S0!�C�)��F۳���E�	����U"qD���D�돴*�{+���#[Y����'}=�%$)��ƫHF7���Z��eM��"9JČ�'v�(@��/�S�Z��Q��� �h���7��XMKë�� �	iJ������L�*��"T���̣�Ɯ@��~��Fq������duf�d�Κ̀��ڕ(��\�T���i����ҏ��ʘ��cb�[J���jD�����8�,�Z>"��:LP�?���Uf����~�o�;*,�8��� ��fΞ���z���ZA�d#��n6v����'-�pdo�xH8b���Q��v��xQ�޺������P��J�@N�w>��y"a���<���1��m�Ԕq�T�����G<�T{M/�'O�MSBSf#�/�ٴ�����Y��8}��]��>>e�7��+�%�P��|<.&��9�aV�����࿧>��iI\��tgV�5�&�������,D�5le�U(hh#��c��c�36��k���鞥D��L]t=��a��S��A��v�O�]_��_��!����|Ow�	)�j�)#�M�O	j�=�r�[�X�M�m����|�@���k���|P"�mTR��ʻR�-�����0'oi�"�D��r�z�+֤�Ohû���E�ehpr�9)�����rnVw��6�r��}�ύ�nSM�?~�^ۛ�����l^f�70�;�<�<��3�J�l[7���@��z���b̫W����4�Zzw���O���r��mL%���@�s,34��2\f�e:�%��3�x�
�>��	�_�5h�2�����"�5� �3t�dd3�Y#�`\�A6�s�F�2�.U
0x7��_0���J�5;N^�]��0�E�d�E���`^�2=JŤq-��`
pL^5��T�7�{��l���g�]k�B���� 蘣�@�Vt��5:�ko�)�R���pwg�u�W��~Os@;-�.~�	�|�t�XH�	â�ΡՏĒ
k:����$�&��	����|G�s)e�ra7��^L]��-�Q���V��ZG��{�h+���Bc�Cz�ժ�tX�(��诧@"IY�����a["L��Y��l��{�)�_�(JM4�ߊ�9�D�F*��b�8u&T杜;��<cdww�#GEsf덂Z��}��;NOEI�(w�6��e�y�7�W.�~�eG�Y*�k�h�^�(�� >5�v="�Z�o����V��h82�o�bu�I����Pm�2	ɭ���װ�/��y�hs8n�*�;�9ʾwԝ,�i��L�s筿��V������w��O4P�{wd�?؞�G��P�h�7�A�	�B'�/}���+|e�#T!���������-1!~aKJ���.P#������azO���na�i���B,�i0J"�B�ȅNr�K�y����V�fi#�]٪����/v�D6���c#�/�J'�O1���Z��I���"z\�
Mt��j�{@��H�����s��p�7�s5���4�4'+K�:�����W�z{���I��V'X@)ﶜ�"0
qzYR�{<�6$ӔqC���]�9R�v�R��{�LZ_!��!�`���I�~0�\�W�c�$��?pR�l�) ��¸�F�s�3�� ��3��l����[� ��Ϊ��q�%�MU�K덙�qز�Ss����0Y�6Q�k��1r|�J&��(�,��D�-I���pf ��3�ځ4&:6�V33�]D+�"�lP�m(�)~f�w��2x}�����cbVK�{+�S�!ZV0��*�4�#T���X�q#Y���sMU���N�(F��o��^�OIb٦h$vN$���@G)T(��X��&�H|������Xr1Y�a�����No�W[���Ll���\�ƶ�t-?];�g�`ǝ͊�䒜�_�@���Tu��1�9�����ϵx�y����]d��  �^ן6^�5cm�q����8� �˨x4]���}#��79s+=@Ť�UD�5	e�f8��ɝ��b���&
�mVd^=��Z45��FV�Ϳ�<&ޑ$���4�����"y����7~jA�����)�Y�{��7h$� ^�~LLQ38�YF���$�4�#5ᬆ�d��ldþ@�P�*.o���k7�2�}Yo����R6�6�	�Io�o3 ��AH2'r�#s�:����"W����{���@�a>]�^�����M�l�eU���2LLq����"�'k�b^���[i퇈��,���|���,Ӫ��%�S �M�c6�Y���O����vt #2;��//�5,UΙ\wnCk������gғ�<*���S̩�S��$x�<B�ᛱ5�<j����7������H���ՠ\�����ԅ��94��,�	���C=�?WLi���4�r�v^Mt;ن��z�#ٓ|��T+ÄA��"�ǒ��>��a�[pg���.Y���������0�R��`:¡yt���٤����E�dC�r兗gNшG���}ȗ3���Uk��s���-l����������
.ğgC�l�XE$Kd'����V��-I�W¤7����//	���2����9Nj�ط�j�z�QN?Ҵ�9X�S0���g%�gA����_(|�[�����F��4��Q8%7�@�mxH~�ѾE,�M����ζ���m����j[�G7Wc�O�s OJ"!�xP�&�PE��G����O�{.T%��O-�������ٸ��cL��f�(2@{W�����@����=����qNĹ-��o�C{�}A�qsd�O�ؕ��u9=Ur&�&O�'�XT��+|r�J|��l��_%S'��T�W#��/��#�H�K���4�{(��J�/�Z7Х1)� ���Yb�Z�$9�� ��a��k�W�z=[�6�+qB.�u�Q'韞m$�����5큮�o:il���/����׫Q���:�o����v��:��_C"���3����Zs�P�vI��{/�r�u�+�D(V�߼�uoni�
��R�#D[x�C�p�˸n�!`��^�b� �Ɛ�����՛b��µo���eН�J&�Jb�^������cg�a�V����q��7hB��l�5����g|6���\r�ڃCY��d4�͙���<q�`��.@�\�J5��~�w�-�%&Ũ�iv���w����9���������R�$��?�L&~����>e2$��'�زʟ��>��c��'����)0#����g$�W,��E��c��#f�-��I��������'���$w�BѨk��4��ލǢI�����7���Qg��ˣ��fgϬ����F|��1H�>���PQ`Bs�%�'��N����߰��L�_B�*J����%k�>�T3&de�㻕l�-�����{y�Z�%kA���KR�1�z���:fP2��x��$�yy"�oQ�dq/c��s��ZdZL��"*N�1�"_ ��\L{��C�xk�ʤr�Q ���w���������`�Eo��g�y'���Ü(�.����
�8l���ElD�]O*Q˵2ڸ��'b��j�g-�pk<4�xIB9��<:�g��HyΔQ��*�3RN�u�'�mLjv�s�.�֦k���K��IG��y��R��l��������(|,	��F���,G�xP�	�ڿ��%Q�<�[ܫMu��������ok
,��M��3�|�1k��7vV�/�8VޒmC�J
��j�5{dJR�k���\LL��<�$���V�+�<S�ΰھ�i�*��U��g+����*�E�"dTnI��2o1<M�$�[l��zI�rw�s�=��+��є�����d���l�����m
Log�1Fr��/��r�K��!8�ؐ@K)Vڇ3o	���P'�LLm�HSU��E����{�A�-p��W*�Ɔ�jL�Xc@�|h��N���4��h���g&��V��H+�x9/g�����.�`Ťd�p��zŌ�16�*����ψ�~�Դ4�'��6����v��<�8D��`?�`��r+�}x���Β����持���Lc'�@E^��"e���+N������VS'�� P�*�J����ƥ8�����;�ݖ`���� ��Cm�S?�#���������`�V	��!����\]�qz��,!l����/� �T$��6�<A�K|b�*�{�\��
R��O{�O|�(yD��[L�]�?����۠�ulV
{�M���9�t
68^,k�	撅���������p�E����Qo�)'w����9����+�y8�n-����U&�ZOx�t~�[�] ����[�"�ఌ?6�2���k�A�I�;y�b�\�I�szZ`ĝ��@������r��Av�4��s[���(�G����Dg�f��ѻ�A��{��k&��=�=�[�3|��x��/�цcTE��h���+}.�[t2�T'>Yp7g5��=�,áb0����r8�J�u�ڐXt��������	o}�1͟d���8��XF5��$����u6�I�0BQ>T2Q��9l�
�u�\秌�	���d��1�ӫ���:�H���x�|��}iT���ѱy�ѱ��tܮ�Ʌ�*���w��E˰��s����~�'�0h �r�_q��6��鐂L1�*���,w�*��˅<fC�D�(k��@O��^&Y�fG5s�����p������� z�#��1���b�a��a�<�������ubu;ݳ��������ɋ�:4~�Bx����T����S)<��>���i&�)I]�u��"��9��*u�\cA����1Z\��i5�]4�u�!�߇>g�g�T�d�{��������L⑛K÷���Ƹ�A����_���?oIJIt���ܘB��)�#�wД4�\">1���P�J�,��gREU]d$Vc�5B���g/>�J��Hsb1�A桇�k��������ɜ�m���#���şs���c#TM�ڶ�nr���We�_!B]n��U�,�|���tG��/?��N�B�%��(��e#�5(�S�f3qŜ?(l�&0(�%?7�����ӧ�a����]D�k%��1.�����5{1vg��N��i��
{GD-ī�<��6h�iۍ� q�i2����Θ�B�3����� 5�{�6�e^Ϛ�xBd���s�.��e!T[��_i�v�0۬�UsL���v�#.�h��W *˫��g�U�<K���R=�\�-h�6`����>-l��^��+C�ދ&�L$�p�o�?Ҵ×*�p,�xJ,A��������������Յ���L����Q�QN�H�F����~8x��f`�Ο�|�'Sc���a �0GP������#�r���/p.�oN̵�|a��y�U��S�o�V<������"�z���d�<S��!A�����`B%�g�t����)�����Fy���ӏhk�׾B��RQ��O'�-�a���W���]U�|s��V�>tn��8%�Fc!�]�������&��KA��B�U�"� 5�A��Fym*݁P�\x�+��9���-��҆լ��t�@0��缝n�vO�T���"D��{$����|`R���'2���U!�ا�/�� ��RA?���ȋh���MC�����c)SlWo���V�)9pmr��L��>��/�B(MU|s��Gj����a$�l"?�Wt�q{��p��.渦�A�s���Xd�X���S��l�-$�����0RWL���_I)�c�E�Mt�.b様���}���%��^��[�5O�fm�n��ȁ?{�+\�W��ܘ7�ͣe2s�����.�ܴKԅ����ԏ4B�1~W��䟕�{�"��;p���e�*D���|B2�����l�Ә�ތ��* dZt��`�MؕN1�$~:L��, 8%o2O��H_P��Vn�@�fj~���q�,yg����8��Z�x�|��J���D�lLh$�6V{���j2��>�Y��Ԡ�[V��Qzrk�7�&ɧ�9�s��C�7lӵLl����uৌVl� �۹��(�W<��k._1�m7�����c��k!�#!�뻟�4�F�3�j�����nWI�(�F��u��+�&��bkX١�} mA����>4���%!�i ]�[ԡ@�e���K�s>����=�Z3���义=�t�IW�@����ahz��% l����D�*�S����R�Y��v� Q�2 �Z2Z��J���蚵P͜��Z:;h��/���?���9
�����=xT��౾�{��d� 8���0�DF-s;l���"b(��p�%<�dxKo^2�OQZF������x��㛇E :�(���V��	I���-/�ϸ��;x��ک� ���jZ�X����� �6�1�A"2�b��
6J���&�z��	����*^��[/� �<�I�/��Х��?����ՙhT��{>J�tJ�l8	�M�Ya���{"���ڞ.��}�]%�g}�_��i�TFQ���j	/���T���
�D�<���v��I�b�Ɩi����H�0]柸���,s�c�Ӿf�Q�U	�84X��j�P�>�K�V�ԋM'i-x�٥���m���6nv�_�
�9s��~�2� ʷ�8�x�r#�{59�U��m~�I�G��i��Y��*,T�My-�S6Mz�z|�cj������!��k�MP+-5�.i��Do���ʭ��v������4-]J#���/~�J�-� ��xD槕Y�\�/����!=z��^�7T������y�٭�ߔ�c�uMm�
�Cs�~���7>�����6�yGg���GW��:�E�tS<*%������[E�x�����_+:_3M���h=5�U�䂼�Ĩ3�܂����Y�5dÈ�Hu��֯� $�0�^m;�GJ���EEGt�l�@�g���}�X�)��Xe�]&�$Z+f�<����|vD"g���^�0Y�~��5$kO�U��� �5����Z��Uq����sa���B�wFg�����ͼ0ÿ�E����� ��"B�R��_,1����fp'3{y�'��;Z��8=���9�䯚q�lA�?Iйm���X�H����'GM$¸�;�(�O�I !��I�Sƛ75�7:�cE�vfz�?�b6��:�=�.T����q1��j"0�e��)C��Y�+��-�]�ns�>WV�؆�LU?}��t��8�1Z�׮��`^']��k!:Y�ﰔ%9%:ϖ#!L�>��˾d�%ౙ}�Ռu
s<F|6�>2�������hm���H҆;P�i�x���e$���ė��ŋ�,?v�Q��h�)�n�}j�@���r��;i&T���E��sE�l;ܼ�c�)�=�ǜ�}m�X��{>@;��;�^�O�-�Z��5�\�y�Y��T��x�ԩ�K�����i?9D���E��Y�R`�4���Wa���b4d?_�i�n��0ϥZB�Up̿��d+�Y&V�
F����&���r�����l.!�٫��r{���⦴��ԉ�v�����8�Rf��q$O�):A(z�*||�5�j W�b�O�qI��Ir�V�OJ�h�U?�T��Ɠܩ�6��<;E�yO����ٌ]0��g�7��3͢�HA�I�ѩR$�f��'>2��.d�	��KY�R�SBR��>��-��tf_����Ö,�I���#���/�����ֶp7$�$�{��������v�?�M;����o��`��H�m�!O�t�<
��:֪�6�K�4�2���>�f��m�6}������]ƀ��= 1k?�2�P`
q���Q������!��a����]oLh|e����s�P������m��M�����z/͉&$�5R��0_�ġ.h�V�Q���%�'�!� ѣ���z�e�l��h.��0�B�8��^�����݅z��?Z.�l���F{�,u�BG��Im���yIT�&tI��l��bmT��zp�dCz��_����� �%ÜE��Y�86���(�?���_�*n<U`�vJ�S�;��i�b)��w-}�H-|��w�^r�������Q�KA�6,�C��󳠩ܖ'�%�T�մ��t��>{옌4AՁO��t>�1qJum{��@ ������n��;�F�ď��d��+/�q�d�v��F�,�H9�o�0�Ѯ�\f�8��?���m�#JH�&���6�C$��8,�<Jg!�+>��ii��$X@2�.'j��t����ߗ�gW�0d�V�H)����w�]L�+���O��\�9�1�§i��7�y�5~�%v�焫5s�^��ds���J#A�Ō���{��U�+Ğ���V�w,:�񬁸�G�b��Nv���=.�qڻʸ����0�sx�N�Hab{�ם,�r��#R��f�B�%U{h灣9�]ӜB�o�t kJ�Ύ��s��G��@�^酈?�Mw��v�2�-��_�ԃ('�c���-�=a+��'��b�K-y;���;����/q>����1s=�k�U{�d:��E(�W%4�n::w�J��1�3�Hk�n��(XZ�\�+?��U5�j�»?G�����v�;�@�Si�,��(�$2o�HF\\FO;&��$N2s����g5)os��?��u��dʁ[�4u��0�='�S��f#}���F�P����[+����ʏl��y��縃f���0�[m�Z��a�Geh)9�W����"ҕZ�U�"��K}zy���(c��$*��ħ-j*˖��޿2d�o:�~t6�����0G W�����%�';���i����"� ��{��u~��Q`?����c��Ak�vMX��_0跈Q����1V����>[�R^�����Rк@�k:�����*(]��F�҆2no�+���R��+υ:f��9_�� ��*d[���Ə��E�Ղ,�����-��~? �W���������F�`'���7lTE��Ql�d0^A�琁#bϱo�r�s�)����_�84In~2���������9���N���I
��zr)�ᣅ���M�����:xz�	���
0
��K�y1P#� IC��[�%�j�b� 2S�nzu���ʾ�_Sc��~��kŎC�u�61S��Q�eG%��4������5E��Ae��Tj���Q�=t��,���i�O�G43F�5�A�>���j��¸�4ʠ�ޣ#�a���z�
����9�+H���;���e�{�'��WA�V�Y=J��L����߳�`���ԙ"�|��Ȇ�i�����l�v%�����8~��nH7���O����;��v���
�{�V/#��SE���6��:BNh'�j��S�a
���3~�U�w<��=�^�^~����AI�S8�ĵ"F(I�p�È�j�N�d-��Xt�G)�6�AW� /��|1�.��T�f�,Y6��}�(��:���V���s��x!İi�Oy���@���-ԍ��7���wH���8h����h4��5x"�5�b|(���=-��S�0�4���*�Y��6X��g���WfUt�:2�"��1[�I�q:iI8�I]f}$��&ٸ$��P��$_��ƛ�3������R������ĥ��1�K�fd��c=Q�9��X�Yɷ���/�`�����RtR�]� �X�\�L��i`��w�ֱFJ�7��e�]�;Ǳ{k�,g;�vR�&pS�"z�=�row[Am�Vq���x��|���%��	s���4P�Iz*y��i���p(�r$���4kN��� �<�^���#��Kx�:Vh���cs���-�Hȣ�t�)00�,�v�%x�4�r��N�2.��(�)O��w��Ŷ̊0��ЇN .ZaL/(:y�ie誾�t�1����Ӈ#�>����A��Μ�w���#�5�b�M��`�@ެ����?��Gư�*|[!'ekD{�2���<yli��5�#F�"Q��1:" ��D�WHO��M�u]@~ �S���}g�}�� /l+��6�É�\�9����y [j�Z�m7$��\������"���t,
q$o|�]�k��[|��d &��p�(���(����0��(M��M&G���U&�Q�'��.�ȹ����ww<���M�c.�׾���6n��z����_[�KUG���v���ԏ*=�1���)y�]�e�Kԅ��&Y�-�ȣ�6Ui���4����<?B'[m����Qc��W�#L[�^���9�|���cUN��.�	��R=���"��b�xB�4�� h-��%z�
ֿZa�
P{q@�ޕ��m%�z�����~�&�!a߂,bv����$�����ߠ��J�UO����T��:cyrmǱ�2�ݏp9���`��]�Ήn9E���;�zvP�hOm���E�΋혷h�T�����Qf�&EM&��W�o��g�b�q���.����gk4R�	��;v�*�y�M,Y��g�m��SC�gd�[� �峴�W]`�q{���Ll<��jf��7תW�n�`k 87��v���Sη�.�e6�����, �S�R��M�����oq�š[�e�f
�Jj�!��n��.�G���**D�pP' �Tc�c�V�E𧶨�f��4��`^���C�a��i���A_3��=M����3��Vl=���_���~3wǊ++�̵��YD�<��	��Y	����a�����n��Z��.��0�5�Z��&�F���p��鑠�xP	n�~1f}���]�v�i^t瀧@t��8݈��:�ܞ�
���huu��Z=��Ύ�GQ_ڠ2_Yc�{B���T���x���7��u�߯j|�ɴ-�!җ��h�ѥ��:��$��'��X������[��?� �b�����D����X��#}����N�]z�~��[6��,�tE��� �z��o�ܴ�%M����!"�b�'�����T�jڔj5@�؄��@��x�#�#��0����L��"�e�"�op��^j�&E&�#�ǫ�4S;�P;�lE4V��J���>gP��\�ETx��Q,\�Ncȏ�,��Ƀl<JN vs�Q�S�~+�y��?M̺x��y2����-L�$���S0Lܚ�P�j��^S}�s��g�|�c�w�q�-2�RǒZ��ݫ�NF�p�k>~�l����Q��<����"���tX��K]i�o��(Ԟ�h�U��\��٧�
f7���tC�&!����b����8��);*��k��W�u�,���y�z�`W�+^0Z �w�e�XXK�m�	ƚ����D��qB1I��i_�����g�q=FW5��#DM���23	�C'�.��(��U�=����c��l3��l��/ܛ�/dD���h07�8�-���cgE��@Nt�3�-��cP|���F�b���O��Ur�[XA�!�q�`���}�+�f��_��=�~ڹ�LQKVqو̠!2-��kvb�P7�������p{dJ/�T"�\.;��b\����-AT�h�מ������|n�'��<Nt�����ӯwϋ�ቦ�$�ӂ���M_���"�R�B�:�Ǌ�H�5�3���r�����K��ْ�nȖP��7e��V�I�5Ь��j�Q��٫&�G#�E���1r켋�G�F6e�.i�����]e��_o�������Iz�D7C]� ��պ5�,[�N������c��0S:Z���CI�w�͠�dd� �I"���Z=�T���1�S��b���PI�_����B�*��.B���Oz��h���/z�c=0���"{*ٯ�h��{�"l_�]�񴂎��Ep�DM�vY�u���h�Dy��:
R��" y�^Ζ�����;*>F�
q��I]3!b"&d&(�)x_1I_"��+���i������6�����o^�O��S<hӥ},+��SaCj-q놠���~!���|�gH�d�� �«-{g���~: k���O~E�kah���+ZIG�k}�����8f+�k7D��Ku��Ֆ�V3��Z;�O3�e<f".��zW돚�����ۊw52nG���НO�a�� �5
��0��n��e�o��"�&�͏S�g]k"̬�_�1M�C��^�&��m�t�C���#�����^��5h���"�j��[ �(���e�^Ƶ.{+�R�T�0��(>p��켇��R7m� 9��4�_̝Фrg'��c��e��䅖�oA�n�m�G��`���N�~�m�X����Q�4�|�U���$�Z���a ���xd��腑�ء�n'L]��N��l�6�U��2REqν�.�jbk�u>�`$5KXm�����G�� �)b��V��
��������^�8"�H�Dro�V�	a���������m��	�$�9
s�ݮk�	�/�'��׀l@��|�J|puk�f��sΪ�2�9�144�@)!�Ţ�hc��;�1oP��[�o��T~N�;΢�%[R$Ȼe�w�L��[�}hL38��\^���X+�y @�ʷ��"�����Z�J��i"�+������"�S&1�$K ��1[���$�g�L0�- �(B���I�FLs ����~_�1��gGR&���jw�����\�{bwԚ��R:�~�D���� ��;��^�@���\w�ᅯ�E4dªy���i�����:�ŗ��J�Ā< 
�b�\�LLN��\ƭS���'w��~f��yaIg�a*�y��PI��y���u�62R�6�|�0��*6� A����j�ۙ���u� ��>"=�����>����B����_1�8q-'�~Hcr�X���Mk~�0u�A���=p�Y�lP
Zǟ.N�Z�R��F���ڴ|�ˀ���CaD������E	Vٖ���n���n���ζ�8���Q@�fR;q�c�Pڧ�߶Q#��#D�]l��L4P��QaM�Pl��M���rc��FȞӰ����sуh���E؋҇g(�c���i/[~0w�t�*��"0��KTS�5�i|�������Ɏ���mpCyo��������H�Zۢ�`崦'32��u���ܴ-܄���S��Nr&��F�pJ5��zb�i �ۓ��y?�U�=)��S���rUXYl��}�����C��CD��D�{�^{����������э��%6���R�ńU~M�ůX,A<l�g�����Q]-�"�Ϣ.�x��	Xv¯!5��
$D�r���Hꦊ������\=@nE5���jr`?�ƭ�~Z��i��)�:����N���-g���#��`U9���-{/�='����	&?�?�&���Bjb�}'f���Y3�H�Y!A���Ã��c5�-�d�Q$Nn�?LB�V#&�`����`�E��OT�w��G��8T"��:;��Dl�0���=�"f�4[�$������m-��1ie��qx��]����߰P�����G�c��θ�)��I�E��ҽ�T2�@�Sa�n��K���9��ψ�p�1��Ê�q������#S���g�C����[zqHi��vk�N&������wT��I�$M̯\?�zN��^yJ�>�9��)־"��/ׄ�^/K"Q��ζ�»�����PF��B�;�K2��S�J��Q��xȜ�S�C%:���_=�Tjx�Ԧ(�Q�Ƿ�8)�	W�.l�Z��Ӎ�#@d��Ɗ�-�''x�3K̟�u��zO���ƫ+�$}�g�T�F��gz�#�ׇ�0�M~E�z���yDb05l�t|+.o�\5�9G���bi�cyO��ޢty��f
ԃ��=�Z����X`vb��÷E&�Hy�#f;�!���صpe����p�%Pr?�d��qMv�x���D�G[�$Z ��;����"up�f����3���/�2��C{s6�hy�,g�>9��R��ft2bp�c\�iOݏ���۰'��r>���)'��[v=� �K͒)~�"^l��G����c��l��#y����D�.|]�\m����.�~`�y��1`#k�=e�0�,7��f@5��z�i�Z�R�w�U"<�H�e�Q�Gh�gu��x#� �;�L�=�RW����]�#}d	��@{kG%@R��1��
��q�����p*��ș+öoF��=�G;9���h�E��[���0S�]w��g��c�VR;��{�Fx\
<R���`K��A���Uu���_�O��
i�C�?�;7�oA/�Io���dֆ�ĸ_S��
���z[tN+��i��'r[<1��6RB�U�M(z_�)h7�4T2 ���)Ĺ��~%��:@&�`.��s�k(������i�TiX��7�]��õ���JI.-憄!�d�'�2"m]2�~0�U��<A���G�z�П�o�?�L]e������V��w��O�`t2l)���oER�0I���G�aP�xK� � ��N���J���#����!E��pߋ���_n!M�ek퉄q	�?�Iؾ�?��4d/B��zh�"��j�9p1�	`4�Х���x�YU��~�<�U+	;_�S#7g��J�HF���j��
�u�r��-jIe5���fw���\��)];��v�4x�����?07݉�B�/~1-���������E��
z��e�������VJ�BM��1�thM�R`�h�F��렝%��|}��b�G�=B��
�{�bc$�M-
ɉ���X�'�/�/,#6�8���� 1�>�%sQ��)�k��9�wD8���-�xXU���h��>A$n��X�-�/��=��
<vͶj�?]N�Y�lC�3ſ~I2m���a0�߁ZI���\��]�,���2�j�B��be$��͡��z7�B%�V0���R��������[�&:C� e}�_F/���9�Y��9147Lj���GQ�5~{R�4�M{'�,?_��9Lm_��^\��v���PiF� �ߙ�*'Dn�2�*Np*i�V�7�rDx�P�~�zp!v�-t ��F�C���Q�IN]�)k�T�>��8V~�P�81�rQ��ҠX�!�-/���p���ur�;Vtp��ٜ%郜�^�^"aa�F ���w���+^�9+ӷ���6wd�M��`�ѐ���Y�*):Ў�ћ�z�Ĩ|J���d�1��L�(DӉ������,�ɟu"�A�,�,��<^L�`�-� vCQ #Q�C-ѷ#��Jl)kd0����#Yh��5���	
~v����G>�z��?j��8	%���K������"Aﱟ�u�/�,"�C�����B��l��)v�n��5�PO���]��f�VZ̵05�x�ݛ��-�|�Q��#w!��Ӂ���kr1N�ȩJ��k��xNvG��Z�	UN�,��3�=��J�*�]������hf�E�9�4n+��bҎz,Me�x�Nb�pe���"3��nǏ��G`p���	1������\�����-w�܃���`�] x�u�+����*7��%0��
�?���#��$�L@��	p��"J����^_��$�W.���c�u��M�w��[�^�;�p����Jk`ht��$���EQ;��<F���:b�	��q}t�}Ӛ�jW�1p>�M�f%�Y��L�AŞt�kH>3x?n��>v�H��������	]����K�	�=�:_E~?2?�I�bc��qI��v2��Cc����/4=f���>H4��dԫnl{�D�K0����S* |�D��̹���J�3���Gnjg<�=�X�',�WW,u7����g��O�ü������,c6��#��f����8;��2�/@HY���CG��W�k�va,jB����z���˔_Q>�W�R�0����uY�F70= q
Y>�ѺL\�.�O�Z��mųR�w&,�&A�_G���Sʇ�hG�����}�˕I����=�8i�W�`!��Q�_���w��/+��N��q@�J}���a0#�K�ϒ�Mu��{�C]%���g&g�tvX��i~���7�/�0!�KN�<���i��d�?:�z�NpZ�G��R<��@>��nW�x~��a�����稴�7��}ǴG�5���]�X��j�B0����*_4('��w�2�G���h:��7%���сٱR���5ak��htyKf1K5�J���I�ӣS�y7V�5�B�0�+���I��b޺�>�v�'�m�����{�?���%��0d����UR�[�{��ًd$8M�S���^(��S�V�񐫩�
d�4�J��^����B���st,�1�S�Z�Ћ��7cp8%�ܥ #9�V��yk	6�覽t�C}�)tn����y�O4�i�+����]9���>�0�f���(�"ك�&�!*��/՜�/�V��$�榌�i7��r��Cg�JR�����_���	�e�MOu ���Z��`�� �󖒲d?�*�X_��>�jR�%땥U��YU�=�P������3]뮐�{4�r�59��
[�����f�1]�rk$��&Y��>�CR�ؐ����w�O�S��J��'�œz� \������܌:6J�tͨ��CF�����؞.@ʾ�	�ɝay�{�t���Q���bE�cRd�֔��--��v'��CQ�0�����H�(�i��㩞M~54`1h�˃�i���
���A�zM0atT���K��s��eB�y�/�k�P��'��ف��P�8*�0pv��i������?kt"����p�Ӯ�\�u�����Y�r��s���f�����[�C���>hM���JQ�u�VZ�z���g��<ֹ8�V�{�݋�9����cy�ΗJ(vʾ�1�(�~�\���0/�4���_�t���M��\]�;L?���Џer������Ke?����d=��?4xt��e�1n��9F�A�<o�<6wڻp9-��"���V�g�,:I?��"��"�wof"*U<�?yE� D�t��
����~�<��l����E��JMW��%�E`��
>�����S��*��oӅ|�/�>+�\n����Zz�P�V�>V޾x�x��-�~7���eΗ]|��$�l��Jgby�4~�r&�Pw��0IOjZ��Ò̞Z�������G����S�8{"�Y��>0�O�W��C�al�wѬ��eL�����5{x�㼢���Rn)�i��n?�u�̇q4 ��e��@b�]�>�T������ P~�,�1lJ�5Z���iW������oNs��]�b�^w�B9��'����ض�>��1�/��3 ��u����dO$��v���s�g���;ޛ- ��W�,>��9��Oޮ��@ E`E&�n�!B��Rk
x��,Vũ�����4���O�6 ���(�/�V�ii�\ c��׶��\��b#��s�.0n�?��	m��[�ݕ��N��;���U����(A�eN���*_x�ITn���>2����#ͧ/^���q�W�D�6ec�P5������J��U-�X��5�W7P�ܕx��~���LlI�ս@}�I������9�ZR�,㹳��dV��[���t��y�f�ń`���n�?W�`���N����:�**�����~
^ج�t5H��R2��Ƶ鎿��~/g4#��q�mq�s6��3�F����p)����Hy��P��d�"��D�K`>2;�����I���[�;���!�p�\��%=�[�4��ۏW����#��
 ���",Eݍ~l0x0���ʜ_���}��f�۞y{Ѝ҄*\s>�j f��Hb�vC���o �z~a��*���W�M�}t0�h>?!���@� ��IƏk,[cR�|ztjB4D��-�IW��k�����dɵ��kr��T3"���g��n�O�d
F��/��pI8�����I�� �S�ӎ����`�&t�&�1��,�z@��8�I��l�!jt�D�!�2�oR�<xU]D(F�o�D��^��d��e�+)$�I�,H���\Ih[�s��H=��g��H"�ts~�����K*�W��M�Ԥ�/7�fI5y�E$�;��JC�D�yӼ��r*���x1�=/Q��9r3��G;6+���y1��B��i�����I�Ǝ�|c=0ceHs#D�y�dFee��!հ�P�_��׺�eE�Aꩿ(����*ݺ�:�Z��.���+`�{cT��t�
%�bO� >���ŭa��z�/�O����s�ǅ�z���!,�<�$���؆RoẨ�mLS9��S8���MMX�|�Ԍ��uUrʶ7X��Xك�^�l�z��}��Z��F�=E*�� 1}�ߔ*
N���J+£�� y��S�ͱ���A<�:���*���8����� /-�,�m����,+��U���پ�T��ȅ��wJw��^�xE�&O�k rdU�D,F�G���D���]�,_4Rc�`���i-d��m��,^E�j��v*�hܚ7x����Ű5�W>�Ҝ��a�����Y��}���^}s| �F����'�V#!6K��'NN��s��X�b��tR��.�^� }��`��ĺ�X}�})�2�x&�ס��L������!�F�~���8�iQ�D��:��+��v�5�����M-�^��[��_L�GN{lg�w���=��=�lq�/���y�,�k�Y ��jA�J0?|Σ�#����`੾��G�Xi����J�re$���{��C����[g�%���_Gs���;���	k;E������)�rl�֌vʦ��B���-�:\��lY�0�&����w7pF��O�^���%��KӮQ�}>15��
)�{���>�v�;7���~H�D�;k�on���z����|7�Ӱ먭���25�^VԳH�`��+(��x�$�9dlPV���^��if�:��N}��_�e�����5�ќ�����OU��0�T��)�kk�ExC�	��m��âj�\rT1I��͆Wz�aA*x[/�W�ۡـ2�B�*����7��y9Yw_����k��5����4���d���0O���{�V~3Ӳ~�+Z��!~�b��2?�Ȩ����v"G7�����",7����.^��B����M�gI�7��a@�reJ��P�3�^�"��<�P$�=�����A���.�y�����|�xR�4��XzMٲ����B�a��i�,���X*8��N�6�ڶ�pj6z;cyG�h�B��?���%me���_X{ٶB|��.ۇ�i��ge���-��p	�TG��M#o�z蒴7��Jtq��������wy��ֲ��t�|�e���r7��(�;TNS}�U�q�fA�6;�*�u���_Yy�{���h`��� �b�8q 7��k��N��1x�.�N|z�RZ�J��U* K+7[��]�r�bl�{L��*��p���R�y�M��6ʣ��4ǟ9y�������Gֿm�(�UD쑀}�G���;��Ɋh�o	˭1�4�ݐ\Ũcܠ֓���D����uq�
��F��*�A��@�++���8(N['�kU�xw�u��{㣤� _��v�0��+�Ѿ�������DB{���Ҳ��̜����؀=��a2�>*�:(r���!�|@��0m�V<��"��>f�fb���*g�Ă�P�d�=Y��נ	�֣�D� ��$�uqu�lf���`�R�S���*Y�i�T(�jǷ[<�t�/q>y5iz��W|�8�"D�W�#Tq�D�HI���&��@L0�F�l_�r�T*�J)k?i�����B�]�n9$iѭ���=���H�:��M�����e��h��ݔ{��k��A�����~�(n'͡���@��j�B����MO=`$�'CP8|d��^.��s���t���Y^(b5)��X&X�A)z T�����ɼ��Oq�p��c������UM%��W�kz}��<�� �j��g<J�$�����Y��U�������zdےyg;lZ�gv˘��Pd�0*C�;*�u�;�b��3�|��p�c���No�M�Ut�7�g/s�,�GA4iY�šM*=`!��-��+Dʂ�����I�G� �ڳr�"�}"&�PH�A�r�FY'M�}�-m.��n��sL��	���>~�y�LM������p�,�v#�y;���d��rJuv�����y����E2�ކ��CIN����]#����Ve������e�D�0qUȕ0�V��L�P|ba$ٜ�OL��, �L���w����?S��mt��Ӭ����v��`J�1�G�A���,%e��o����)|:��5c4Yx���߲�;�,ި&:ɩ>���q�N��
�)��| �M��%�{8A�� �z�\~�W�Z���A�����(�1�����/�V����[������̺j1��πw,d��۳&��Iҏ�0��Z잋-
�F�Hy����7���p�2{���
ߩC�[ˋ(��:y*�.<-ց��톀��3����4� �m���ķ^5@E���q��*�I����$tm���}~s"��F�aVp��ޠ}W>�)CB�0KЄ�yƕ��<���$#p�M����	O�B;*�v�;SSq؍�����j
p�5��y*!��iMJ<��v�[�S/)r�'GD���Eר,)C�hU��$��pl��0'펃�ƾ�&� �qi5�8�l��W�7U��X���z�\�&����~<v��]�"�y4�2膊,|�~���H Z8Y����қ��?~��S4�� D:��C��P��d�rB�5��	7�M�n�9<��p�RG��h#h��rU�	D�pwG��d�O:@�@3�ϭ�k�l�46���9�%�$0�R�<kc!���h� 1Kw2�l���͆J��V_11���� q���|8"�\���g�$�O�nv�8���T2@w���; E*��A�������Z��}���DdM�&Ɋ�D�֋�:��o���Bϳ/ٞbTn^h/��8��Ӗ*�<�T��*/�C�(i%�#\/l�^��5�N�n[z�ᝆDUf��<���q^��h��X-晱\�e�a۵���k{D_����[�ǡ����K�7�����eh�I� c5f٣��)w��:	�3 x��`��A`�Q  _Z ¥�ob P�|�e�$�s]��K/d6���xO�l<�2�1���$�:�
>(�Mq{�P�4�5Z�GE����%�Ư�u*ԣ�HIr����2�D	������r��;rm��iΊ�UX���ϟ,�]�)�;�@�.���j,j:��I_�G�=awCd�|�D��w������Fh�
��t{h&�?�.N�0��&�K�m���X�x{
��<��·�?B�BTm�=�	_�򳋒�Cu9)�����q]���g[�6��p�ݼ�R5*U[��&��u3�^\�*��' ��j����c��]W��LB� I(_���qm���_�W���E)��_ض_�떝�?$(��(<x�^��W�%)o���E��yy��ȷ'�o�I�а�@��G�'W:��ⷾ�Y��E]6��b�+i�`�w&h�j���U���~3�d{�+s����DZ�G
�oB��juqbehIM(��^����X�)I{��j�`]���|^A�:�=6���9��`�z�bUVco�E:�=��5�8'KT��
�3�8��4�BQ*��xt�L�1;C���͗���C��3���Z;3�*4�e�睩Q��od�sx�h�M���$k*?O1���O��jE��;!z���{$�to~`Ed�1���Ʋ���*���_� 8�r!k��TڎIl��M1�-����GC{�΁����}�l�
� ~���F��U�2.�ɯɆ
.t�*Ԫ��X���	(�E~!�X��'^�bW��2��
�X�/HV3:񺔧�{G���0Ƞ�k6\؆y�}-��Qb=\8�/��N��S��&㝆f���{����a��v#a��o���6�۫Gb�~��kyT��(�ÀҐ	Vz$ASe�3I�,���i����ɒ�ۚ�����sg#�ݫ|<OJ���v>y��0��8�j�8&ѓ�	��%���hg|w2���厴�|W�9�|y�&Q܂i@Nt�|�wLl0��q�~V&�Z���p��^� ��$���oR##��=o�9���`L��Baz��r*���!	��ADg1�La =کy9x Q~f�D����L��Rm�C5r ē�Ƃ���t��B�k��VKUG�>6���kD�+��)ك�$�K ��h�����t3A�e�tQo�s���Z�$�������H�p�tՀq"�vp�������G����A�Z����՝J7c	� �	b���&���'&��m�x���/��g�:V#�jZ�d���	>�11��WO� o*d'�Պ.�����g-x���B�S4g�	��x~���ĜH� 5��krώ,V��E����{d1,�j�ny	��Hҟcw����߮`�ۭi^.&_�r�ESd�~c�Qc4�v���(y�/�,$A�D����_~�^m���o���W��~,�$/$�I�OzǱ�Mt�~�N������CO�@�a1e��=|_r8W q�Zb4��j"H.c�f��葚l��G-�/�x}��"�(V� �}��?�P�XQ�71`�g=#����8M��M�e(��MrKVGdHʠe\�rt�99
���q?�O�G(8[�
��;�����H���SY��������^៊�	����5��}�7$�9�_�;z"@ooB?��߁�,��L��޺�9�H�g��L�$�����cz�g�ߡ��ҚG? �E��v������SشU�=O ���.��F$���^˨Ln�������wR���$�W~r7���*f<l����H�T�OC71�W�ȧ)�͉2�=#��@�x��#=Pd��eP�d_�nFȇ6*_6����৮
�n���t�5�a=�Mx����{��a��t��7lD*��uye5рi��v��4"���,�)u	�o<�D�Ǚ��Ŏi
m��my�*��a�h�Ģ��iW<Ae\�&���IJ:J�T��I�Ə�}���f$D��_<�Bn.,�٤�٬�Z��I�?�����T���	�z~�89��FM���쀕2
�o����t~j���.��-}�����O\���?�Qݠ�(ԝ�U�l�jٚ�-	OoM�����R#��LߎY�̗Q;o��ؙ��:�����9�yۖ�����Z�x.����f��ǒ[FG�NM���B�o/�!�S�V*�I�k�@	Z"��L|
�34k�$����M��%��<����1�(GV6 ��Vև��y�Oȷ��pɭ�#�P�"�Rx����x��Cmc9h�ʳh=�*�c���j tL�*� ,j�x��R���K �\A����"���h��
z��i�g��p)ךó�)x���7gYNI��5J��#��e9"*�G��+� �Gw��tMn�7��R��u��Ĵ��L���Y�J��o�i��u�odn�!⿍�������Ƞ���мܻ����n���pd�=9�m��Q�p�u�ea�a�`ڬD���Q�������R��4׳_r܃?��,��ް�+�O�F�8XC5Wդy��DR7)�2P[ �uf{�馲7�y�b����A�a�KK�.��m��Y�Σ@c|��|�L��s�[륥���՞&�����h�yV��N�̼F�Xx�%$_��)��Q�5B�㉗�Nk�L���c���_�gGl�On�Ȋ,G&��ir��c�mS �=�*�U0� �3�ɧ�dJ�]S!.���)�H���?ɗAjk�n(���3�Հ8;�~�s�TZY�����+�,Վ��7�[��uz�R
�DkD��Z�j�RH9��?��7%T�c����q�%�Z-�_��|�X8|�R.r���)���nc�w�}e+/6k�C���ʎ�z\ڧPq�H�mԾ%�a#@���f��R�5_@Jh^P(��>.�o Ή���b���s��^3�SJ�H�)��� �'���X�N�]Qyeb����	�ý�4'���(�T����@^=�2P��	�1C�&��ۜ.h�8Z�"ɞ�\�u�\7�����X�A�cGC�n�m�F.	'��8b��膞+ ��˨�����X�L1wt�)�̅E$��/_.�4J���A�6���y.���n$$�v���%�%��8iO'b���#���c��P�)Dip̆V�^� D��9k��V����-���J˞=!N	���KɻTj�/��H�Qk�y����/l:�Qp�ȏk'��17����p�]|��s�[R�,� cL�p�2;S�C*�� "����ucŇ�R.Re����\��`����R>Pޭ���h���t�~ѷ��L;"��y�ԭ;[���)���tB]M�+����A-bM�_��r���Μ��TX��Ԁ-�q�Av� M�d��X;�iGb�i�|b��}�i&��"�o�L>�������� ��96@{n7ܫ;���̶-:�%w�	e�;�Um�UGZ1������;@��2���J���|����ш�q�s@�E_�rw�|e%;�A�;��QW ��5������ۜ3�����B��;Pa�����<O�_��v!�18_�
­o-6w� ���OY�e�~�H���u
��
�6�<�Ǽ��x��n��[G87'�\�lu��ϔlY��=�ظj%�D��MU �C�=8��z�	�DT
��Cޛ��e�E���2u"��1�cg$v�Wz����.�n���@�9�7�Ք��4n&?q�6��7SJ����-�~'��G�tp��}�O�ډ6�"1�z&�r�9���[I��P��Ċe�};>�ݭm�I���Rv���d�ȣ|�{�l�Kq��ED�b� 5�2F�����7"�-���J�F�龵��-Aհ�T�؏9���zX������}�^|�'�����W����,d�Nğ�"�:��{*���Ɣ�,�4���(�P�L�c�o�[jy\�:>�:��Z��[];���Vw1�]�x��p
����x=h�kqa�'�n�{�S�T�Y �6N��w�5sw���
�����ལG�V���]����pnCn�j�v��x
Έ�5(ϸV����@�KjH�	V^�X�t5��G��z� �}����Ki��U��y1���(aL�cm3��B���\Ka�8��Y ��uN
Z��&��/	Q�%�
o̿���A�p��U�{QDu̢�*�\��g�J��O�rŅ@@��3�4.���b����@�X"?���E>qU�M���X,j�u˓���P,$����ɠ�Fg�A�LP��O>3�mӧ]��U��5}H-��1#�����a+�w3�;7f@m}���F7�ku�A��x���:�B#����t�,_�,z�2���[���k
�r�%�����诖:X��ܽ|���y�)P��Nq�_����39<^ڛ�cY=���M�w��Z����+���`}86�~�i� Ut�P"�Ù�8�PeG�`sxS�m-3])��T�#"	��Ʉ�cjS*�U�����˄�[�������d?}c?F\�y�ak�����g����(��W3}ҟju�Q԰bd�g��UENv��t�c~���g�Llc�1� >y�cD���!V���I}��_<�#�D������n�6�����Ч'��H���U`�H��:��W��	x�b�z�}Epb�����;C�ᤴ�wss����o���Mv���qff7U=IUh�2s.U]G9�.��0_R��ґb�?n ��F����2bb/�5FS�h�Z���;�h74G���~,Z�O0���D��M�q���������!�v�
	^z�L�U}oN�e����Pʬ���'5y�p���<��Q{��W�I�Y���'	k(Y!!v���:٠I$�rq�&�A�*�K�80��XZ�*�u�'�''/[˕(�Yi���׳{���4"t:G�R���X��(��t���|��/8o�4}]����4����><���+3>l��}�|!0i�a_���ޒtN�4�d ����o�ϖ-q��2\��P�E����	8}�����v�@x�,
η�k����Lޞo�w�n��&�����pv$�,'c�a�F�������$ؙxt�x�rf	�!��8&XxO��N3P������Ӗ�sf�&���izX�"v����{3UhJG�Hb�`����:89��3bҭ��^
(�m� ;è�xQ���͟K�Ez����/��,H���[��ĩz���"�*�I����P���*�d�bH7��>3*Σ�+I"��;���޺S.���/W�g��u��0W�T��,��	�����w�:]:��6�cg�o6ɂ���c�<}��J4 w�E�cC�}�ںg�6�W@��(j�ʖ��јNwtb
<`�<T�B��Ghx�(p� �^|�j�־Y�5)�Q��,����8�Z��|��cm��(��r�uoW�_����*=~���z�F�K��{QH/PDi�����k/���G�NX���z���6�H�R�jX�ȡ�����Q��w�g����^��8s�O���V�nto9�`Q��d��W��[�D���o�H�Vu�TML�"��MS3�$	е�&tBG��������M��A�z��`�϶n�6�X(\Ok����Y���5��R́��^m�2 N)��AI��R	85�ꜹ&e�lWn��t*�P+���p'�{Ztrx�v�F��몢c;����#�{�Fߒ����=Ĵ�j�S��v����|�;$X�jZ�&�.�{�zpL�`�E� D� ���y��l�:<i�k����8}7�c^P�_L�(�|#�gH��5����i��y��Lu�V%����vh�
�	�@�_xA���\WC���X��L�OG�e���ڭ��#��:��=��9�t�~�0h���x}/�������a�ޜ��t�By&�]��}u#�o^��B�����h��Q0�R(a��%�n�jn��<���P>#�U������>��j�]FR�d����~WN���:��o���ŏ�v��.е����SB���O��~IhlI�9��8�5��Y�P��7���h0�� �ؕ�-���'���{uU�O���R��ˌ'<GR��<)�s���E��C��n�}|೶���`_a�>�鶌1��l���v��	��N�xD�3�9���wU�+����v�����հ��U˅�r�z��֮�W�d��X���}���� ����h^hU�'d���+����n�� L�!Bؘ�L���oGY^,�פld�Tz� ��W-˺p�#�%U�+)�*yKE��8Ǒ����-��FHV�$�bL|Ǹ�W{7�����e��E��E��7-Z�k^�n�_8d�������3R����m��6�E���a�e�Fb�neV��,ޮr��E?���ݍ�����i�bM��l��+0j~ n�Д�b���f��q�Y �Xv.�p+IWQ,OR���(o?^���Q��h�nTq������ˇT̂_����-sE��%���8O�
�<kE�\�f�����5����d�|(�bN���UZ7�Ṧ�t8s�#�聴�V�L�#�����y�ҷ�̵�&u-vĸ���l]e��+@ `o��}�

�P�y��d��DF^�m+eÿ<.b��n�q�s���E2ߋ?��%��,L�B�}شO�<��a�!�k8���$b�z���]��J\�E �
�$nfG�aW_�n�o5@�+T}Z�;DQ"��"&ps�*��P7��>LA�p&�rcW���qV����E�$	�[<g�K{�=�+鳲c!7}��F^�v��b��m57�gj����ؠ��Hn퓋s���/��1}�'�X�<Ď�w{Y��σ�b��!]밸g��K*ƌbѤ�Q��+�AC�gZt;�y�=u)����od�`�x6�B#��am�M�N�Jh�d!ދ�$�{[b�Ǵ���q�˵f,��ç�	�C��d��M��%�um2\OGOȕS�]R&ٺ]V{[	�~�YGh�7�@��¹^H��,%��&_�-w�aUx�5_�}���C��+4�W0k���?x�L��r��2����|��ъ�X(�1
V���r���b��"C�8�)+:��䙨J��Kg۾�v
�z�������h@�E�)�I$��L���_�wa�)�w�g�ゼ��w��,�f̃�&6�u�h�i��N)�g��.�r��+�!���f{�_�7DX^��csっ$�!l��l�@�ceTʿ�0�J[U�Hp����
Э�oo�c�����i=�Q��M~�/>�t��V7]hb������;��4x6���NzN�sY5���F]�v]g�*7�/D��+��h �r�U��#���|�٘-h\*�H -�S�����6�t�xa콞b�\���`b��sT8���fx��~�E��;�?R|�Ή�zJ���'����V��3�<�HЌ{hq�V{�j6�%a0D��+�䀛�7&,�8����e��s��X����%މ�`i}˸�r���"�����t.A����ͦQ/j)���_7~��%��}h�2Y����� bj�����_�[�*q>����2�=g���p�[�E��s�x�ʋ;K�X%{s��5M#�h%�'nA�� jlax��^g�����ק4�&s�&9�D���݉4%�u�tCY#�s$�������3C��ߖ���p�Ѓ��|Y����G��q�O`�|kwҁ��v��Z�Gڋ�C(�X2Na&%%�];V]^��k�+~��ʣv�<��5�8ᖥ�KX�j�ay�A"�G�on�q�����zHǻQ��/�͗�o���Ǌ��s"��`�cĆ�w�IJ"��e�a1�d�)K����&}��ѥd:o��_� f�c������2ۏ�&
k����� 8��B�v�Q�I��6~��A� * ���Ҁ�[L�V�i%D��P��z]0��N����yr+���'�q�O�^���I�d���CWGW.B"�08�.���ٸW�W�e  ��T�u �v~PsV��B�V�;/�ދ�gs���S��wiŹ�
a��i��V"g��ޣ���/������ѩ�2Q��cܣ��s&��CfR�>ߞ��v�tu �3$����y��|�k����d�"���{�z��m}W)�w�L�-\8W���%�J�~{h��'�sǟm��r��b{^4���ZR����	v�z4 �ۛl��ō�gF�T� ��)����o��iz0^�U�2�I��]�+��.�U����
����:ei�ms�l�x��ϲ�fSuH��b��_sF�5x��S˗���:�иu��.�2�]cšV������?�ZZ���>�*�f��'y���Lޢ"���м������})QuĀ�\��;��y�"+�K���M<�H�N�v5n�r(<[xH�rl�^�e�z�i�^�����k��t"P!o3*i�Lq�\s�HCw�< ���o�I����U*1� Zg��R�F_{H��RE�Fϳ~>߃�Q�o+;L��^�9��D��pJ�����OV��Zj֬#���*�!��������k��@zy����1E�J@O<��U���C;.��h�}l�Mۢ�H�<��'�K�r�C%l`u2�i���'&=�/�%@�u�G�c��/4J��1@�d̩����Z�.�����Z�
1���~DFS�i����ZP+����6��>m�g���
ט��6r�X��Ǔ�L$bFuY,D�ݔ��#lwT�J�'�lUP ~_�o��/.�a�U=RPii��3ZA?I�B)&���c�.9�LJư����d.u�(/���-J��"Z7ֹ�o*�ɫ�t����zC����T�ly�Ӌ����ϙ�k�����76�0K��j��0���f��&2u3@ʓ��{��Y>7��ü��'+8���	W�S��ˍw"X�Q�����,�B�?�[�J0�|r�� E4���ޥ�
0>4��*12d��$���:o�����)��TW��N�9��z�sF����̏����>��C�9.\HOڲ���,[2Ȏ��{��/m(t�<}�{���A�+@HЃ��y�W
X��l3��ue�p8^:Â��CF>7vm0��nw��Ex��3?�s|}�bY��fu�pf�����f���\� ����o�7�=�0�R����� ����W[,�,댐���<+[	��_lH�������4�	\��\9� ���dӻ���MZ:�J��C+h	DG���7$�ƹ@T+�CH�{��I�r���Ef`�ҩ[��"�e�1�rӤ?��ٔ�3u���*��Z)~$%`�9����!����q� G����Pj���8���-�x�^#�-���o����mo�t��޷�	��Fyv��@�1�̓P���h�%M����h����Yq���l>�C�6��Ԭ�g�� (д���RL�!tR�I����p��ѭ�k�kY"�t�n���W�z��]b� A���J2�g�b��D��4�B�JN��K�%�8���`����"�hv�9�o@ �����/�_�G�;���-�^��V��.z�a�A�x[�o�2�׭gr������>�HK�����6�qQ�nB�DCwa��fy!rH�"U���g+�P�ו3�uh�bwDoTו�-5����o<~�Z)h�ΰ-��u;��S���s�g�^W�*�N�oU�21�#��uQ�͆Ʋ1���$�Ss�|��Rb��T"�X�Ikө�E��B! �`>��߈��NIP�s�VO�Y����u����^�y��5�I>�!��1�M�Q	B� � ��
��cF%��9�v%7�W6Wլ@?\��*�8}���yÞC%p�^�^��WCP]��*Ž�݋���E�e7��a^��'�MTN�/QZ%9H	���l�3�Q�غ�<�v$.�АM<"���@Cy��*v���қP�@P������P6)��5��UUo&&P�����	���N7���b8|�6!�i���8F�%���]��D���xN��[��࠯j�h@AsP�]��w�<����)�+Y*�RS�pCha�MRL��@Ϡ�čn&2o�,N��j	�_iT^�m������2l�+]�s��9���¿樢tp�����h��@>��zf��@n�-}4�-��Bk�wk��ez:Ď���֡e��Yi	9�*�����표��>�A�*��qu+�p��a#P���b�"TR�cd7�[:|ѮZ��
���8>t���~�v6��uur��W����|,d��Em��|OH�x���J�z�EQ�4�.�ȓUh ��N�(Q�?�0�5G~`�4�<�[�e��ӝ�m��2���e,�y(��#CVh��ş��'W�J�O#*��Ű��D^Ļ͇�n�g�+�q6)P@>	r��a?v�(%��pKX�넜^o��Nd��H��Q��P��� �4���KOq��w�g
�F��U�U֮iI>�nv9��q�h�����l��¸�:l/=�B��;�<�'��1{RN�l�q�w]Օ��x3��b��{�-]���c�ƻ��[�z�_���I.�ް�(�ȮGx�c���k�N �$�;�O&�<2�g����Q}�`��I���/��:�?]�SH��7�Զ�M�Ȓ�� �߱b�N���(�[xq ���!��C�����I����3�A��r������I���m�~R��m����<�d��uKE�HCݝ�L��������2�}J� h�mZ�y�B[Jo�SL/�)r���	*O���U�j�w�`�W�A��AصQ#�D���?�Cm�
��f&"�7fkSB3����W:o�$�ƻ7�	��Vy����í�T��A'�f�XÉu ���W͊w���<�ݏb�+�ckY�M[�m���g8�+�\��v��I�Vn�J;�-d�]eL�����}�����c�5E�tϸxS�u�}T����>|���?�0&���c���y���2l�2�f���?���I1*�*����/�I^���t�I��l`��^ۦ��,Nn ��-V�� T��Bυ��|� $�e�9��N�_/!�.vܪ{ү8�Ib�`~_��B1�2�G���q�28KO�q�O���*J��\M��3�ВL���5�A�<�r����#�$��P�bqSS� �sg{(���}�(� M�ː��Z3CS��S���q:�ɀ?<qRj���<ހD��F�D���.�X2��5"�$�/Խn`��� a�?��{9>>�+=߰O�<Mjz���&Op��5��Y ���o�1 ���[��<3��\(��b� =6|�:.c����.e�|�f�GJN���˳~jI�ǚ�v;L���j6���@���ȭ�ădcEr�q�Ў��cE��s�-�-'�z�<�!jܜ�������E)�*=�N�D��{o�c��	�re�4��,��ma7*���~R��Й!��P�(�V����̄��d��ӑټ�wӦl:��o����26�}ԟ��|���>͠��k����P.^�N��Z��AR�e �c��*����0zG���@�����F�B�������K-
gY�c�~;����D.�?��+�L4#�U�nE��V.�u{C��0�Vֹ���/����{R��A�d�IǞ{a(VG��d�Dʚ�Z�o�G��ʶ�$�� � a���*��D�B��W	���݅3,3(��D�$� ���K�&����<���<�V���g7EowT�����"�����_�W�7��؎P���H��Zg̖�J)-�v��_�.q��MUSb^��*�p�N�ȡ:�b3i����֏��.iLb߱u0=��w�;O��V�2w��"�E�����X��5�O�Nk,#	�Ad���|c~ꂄ�.�/~0�Ev�L>��{y/\�����J���c�a�'�((��ߤ<Ʈ��.����cꞋRO� �6][�Oy�r�E�th@Y<��ʒu*������W�Z��,��̶غ�yW$��I<��XT���Q��3�.�oF"����P���ٲ��6_���w-�6��Ֆh����[~Ů�q���+�Ҥ��2Y�	jC.o��F�-& ��z��_oPo��D6�����B�b�9���C�2��#��R�*%�>�d���w4���2jt��Ѻ��6�%r�Q_r��RAP�M1d���MI�|"����g�mV�p�7�hp���K�X&m� ��З͡�m_������
��Ew�q�.�ߡ�L�o�_]З�l��ٰ��gxʝ�4�G�擤��>�2#��I��
����BPX1�ٙ���ˇ	�ؑ�ጠ�5�yS5D��ސHV�P&t*��!K~���Y���q�X`�;�Ėz9�V=e����JK�I�)��Гa�6�(��2��V9��[�+XTS�,U�J��q;��WH��7����loM׷yCԸ ���5��ʞ;��\�2���E�U���&Xp��~��T��d� �b�%�kT���������T�^���F��& ������>��Gq�4�m� k�2��������2����4u�@�m��|'�b�t��(GUS�C���������Y��
�&�u�}"��v��jv��|�u�2��#�s��oV#�������tL�i�m_n�.B
�B� 6�>	���$�'TUNgEۗW`m6� ����O�z�!�����)�T0̓��?�V��4�y$ON��������YAh�C�v4�4q֎��/���)�����`����`�#w��(�5&�-�.����&��7���M���ܖ["�	�"V�O�6�L�(ҭqiл�B�:UrA��wUV5�"����h�fb
�A3�vC�n�~&���/ț+��,��c�:}���ߧ�\`�e�:��l9V{$���mID���n��l �|���H�88F�Xz z�Φ4�.+�Hq7i��xSq�����6q��`�]V�4��2��������E��#k��&��U�B7�����i<��������w̃g���j(��Dr<n��gi�rA�\�?�����N�ӗ @�Y�ʔr���q����ژZs�*'�<@V8��u�?�_���
8d�⡾CC�h(�2L�zS�Z�؀#6��? .�NWqd����,��C�V�"��7�?2 \C���R��h|
=h��7JJa�_* !���m�c0Mp'Dy�~���! D���X)���ʹ9���n���`�(�j@���@�8w�/��w���7�I�z�S����-��XB3�/�u`���a?�*����S�+{/���j24�VE�<�3��0��K��u	P�jծU- �|�?;�f
�HN�r~�u�,ݢ�1iAdϸp�`7�1V�CKo>cp;���Jy�,�6<!�\W�ͫ�[��mp&���#�&�V{���j+�b
�Bc�PY��j��7��%;J{9��D3�G)M��}�	��v|#�D����ܘ$j�������"���KK%�o��^{��)%l��yG��q��yJ�]
��!ԟ����}Fy\��!f�.9��G5y�Ʌ�!�>��[��y@�O%%�~�)�9���-��M-�X\y��l^ܯVM�����S ��~�2�k.��'��i��Z}�7Ji�	��󬽴�D��0�� +Ѣ.P	k��d��}s.@B ����C�}�+I�9n�Y�����~w_3R�ɗ�Q^ws�9^f\���v��uH(<ZN��.���Ym�\`p���$�,�5|��2[�NX������N?�)-6aI�$l$.yE��s�0!������"J��V�&�	����4�Q�wa���M��o�U#dO��8�'��a�p`8*	�Q��%�|����Q}\�>Jh�p���j�iG����?
N`�717�&M����o��0�X	g����BQp��J�h��3̦Ȫ;��.v̄+����L�;_���c���Y�X�!���<S$@f�)Seɶ
��r�B&W�C٠��ĺp�L�6R�:Q�;��X��%ǥ�Z�����3m��@�[B3|&v�֬Ǜ#ږ�L	�)	J���H�,�@d�	���� k>�BC��QxՈ@���*�������I�َ2�eޢPj'�aY��!y������z��u��A�)x�\�r����b��.ށ���?��1ұ���q����
�����[��u-�; R��Q|����Íf�c��t����� ���+Hbp-�� }[����/��@�w��D�'�V��3��5�;��o�&2�A��a�E�$����v��0.��:=5���>�
Q������6�� ۟uiT=7�t]��ao�"�	�~)�"G���Z��M
��s԰��k�B��4	ʳ��!�.'��
��b�aY�1B��N�4���};�#��V�K�z�=����\�
A�N]�E��{�6�&c���r,�u��x;�X`W���ЦAa��9E�)��8�\	_���?Ə��t\�ٶ���Ls�����ޒ�[RԢ��
ߑ'�5/��~�ɜ��8�zi��V�D�}��|��(A���D�V �h(nh���W/��_z?LR ��&�����в=%hXxC��LQ�:#��Go���E���X�a����x�z/3R'�:�ΐ-���dOg{�BIl	���@�>`��؏�9_��F�����"����-�z��3c�˯�J
��igk�V�hs6����^/eH^L��ݭ�/��c|�y�i���,FLe���Uj>�/���f1w���@$TQI�_y���*�K�L �tn� L��	�_�?���.��P�Ut��9߂Oq^L���D���9W�K>xY��(���`��SW޼Ca����}C��EA��L�8N����,/�NAe2

+�F�搙���3�@A��Nh��jo��bUS1+Ar��@��h1��2d�Dr�����U̢.>G-l�8O�kǟb>z����`����b3����J��#c��ݥ*��!����nsn+1��]�*?$o�@�W�ur]�rwY����T�s�sA�ڎ�䩄�t8����%�<(o!ސح�|�3�,���6?�$�0�4�<ȯ^OEr&��W�|�Ż1^������K4J�{��ෂS�+o6���^��DT��g�ʡ 8���@���A�,!Ƿ'��d�s��zӡ�ؘo�nA���AY{T�9�})Uo�J]��X>��oܘ������k��q�֥�%���t�3Ю�D�;��pΦ�i��b
aQ{����5��7hҳc}�fG��5�H���V'H�dF�s3Y����Փ	�%J���O�'aY4ǺD�6�H�iT~�����hQ�S*�� W�]Q_ ���%�mR7n�{�O%��K$z�H����-���3[�_2��v���=f	tf�7&�Y��,➽���ϻ6�Vq�G�xζ�Y��'�����ȩ:�F#�YP������=yUnA�d�Ռ� ��i�����D-��j�4����?�ܲf��ո�)_~��b��1��Up��j�� �S,�,��5���&b2�Fik|"z��Q��*��m�v�+U�f�#�rm��]o��bl�����ٷ����0wڇ�9�x,N4�i	��A�yYrD��-�m�Y���o§�f�+�JC#����B����R5��F�+���Ho�M��?�mq����C�X�ܵV�\�\X�Ѡޣu�҇��ϕ�4,�:�*�^E:�ȫD[����Y���5,��Gh���5�2��i�D�@�C73"I�Wt���e���=ד��	r{班�%��\��n>�o)�T�� U�:�1�0dᢡZ��}(*�T�:��g�)�jH��A�_c��c����Z����c�`ldn�L�I?3�[��MC'�C�Jқ�#3rmRWQ�(�2��絡e���&i�V ��E�W���z�By���Ŗ�wUݣJ`�7ޚ`x��$Ms���'��.�X<�����L��rA�B�v��8������� /ZJ%|�V���b�Ex8�b�S��|R�i+ef�"��ga�ȉլ�e����SO��X�ڽ�����/7�sv�+�d�؋�͏㢂fC�F��M���Quj�_��$��	��g�M�!���RTq��Y�G^0}�*�o@����+��f�"`{�{!�C��Ω4{��d
��+CkE7Y��ߘ�h�'�.x�i6�dPW+��K��f�w}�' �Y�)%�[9d:�4z`����b,��`�0K"�l1�'�u$B
�#��v��=:R�5ؗ��t�0�hC���������&��0�3�Z�wo��!������6A�*poE��$v�M��!�6243�6���Z�l�Uyfo��*J���^�ͯ<�元X�;zٻ�}wK���J�B�|R`>�᧔<`1�?6�������Y��;8�!;-�}�F�|e�5qGJ4��c����u���?h�K�5��&�F8G�A�>�-� ��61�^;ń	�����&��}�;a���G#o��A���@\���W�U�$���՞�P�d��D�cD�9���l/��02Cd�0/n��:���ߧ��_Dt9�D��L]���Q��U��<��L�g���?���MLR~Z�lcua�qJ�ַ�L�Q�n��4Ki ��-�ra{³l?�ҏ<�&�z�Apl�� n�U"�nj�bMF�
����)
N?�F��}2� )F�TR�yX�&O8b!sj�^ou��-F���ln?��U�.А��VqG'���W8I�]a��[�	x��[ 2�E�l����8�$�<�RU2|Y2���IK��l@������1<�� :��;=+��φv'�9'���-35䘪��P�p|���o7'g �!+��ޡ���ŵ���w��R��h�!��8�B� �ϥU0X!o�L�����}P�|�-�
%`%n0ć��S�nQ$���_��zĂlY�D�ފ&%���"KG���)�c�T>RF�x���(.|e	(��TH/��K��olq-��� �6}�Ԡt9"pK�i�;����ȕ��vV1�e�W��τ՗��'��[����!�i$���s�t?|��P�N�9dc�ˢ���raЦ\)\�|w�,��gj�+���R�}]���H���J~�i�ե>����O4-Ԓ����d�Wb�A�����ǎ�ĳ[�ҧn�-=�=���BQ`-+��oYb�Lu $���-h[�������w�_��A�xQ��3�M�T�H�x=���&�@��n�ô�d���8~�k�V�a�����
1"�����Iew��/i�e��2��m��%����h1��w�kV��EDW') Y��Q_ G�yg���f�?Qn-�ʖ�	�_h�Hi��ξbIU��:o�U��l��tD� )�Grs�*3O}Ә;��U4�\�0� �c�u�%�8S���<I�����XL�e�'��,�QQz���򗃠^��P'�3��q����$^<u*t[�,6D,�X��[�j���~��&��Q�F4'B�'�ۏЦ5,��%��_d�\�Ցk�>Xybzz���x���n~�O�k_�v]4�Q'��\ƠչA�`�j�����'���ͳ;����ʩ���{��N�=zmz��U���c��d�X��~d�������%O\7
D�zN�%r�@��Ӝ��Mj��ڦ��ZvX�D��]�8���v�����Q��C-��#d.�������wz_�,����<-5�W|�җ�]�ܡI&�hr����/i�\$}l��"��B�y���2��8Qh�W�}�o"\��f��C<:0�������5[��M63�r�)�P.�oi��0�+�抁-��+��u���j`[��9�$���D�r3��}�F�#�zS�mS4�w�Mq4K�y�.q�s�>���i �ʣqX���b�������]D��H}���gG��tk#����
�!���^v�1�_M��:~����h�_���p�+���
r@��o�b���舏"��&D9�^��G=Oe�}s۩b�!s� ١�r�I�^�2���@}�l�7�t^�;�9�G�j?ч��
�Ӡ�k�B�����p�_r ��#�_��=0��2�����/���u�?��?��"���
^�5��@ˈ�ݐ!�h"a��Y�I����� �$̥,*J�Y5߬���wU`����=ṟBi=r]�e��~�mZ��$D����`�l]�o��zfh�VMl'|Og�fX!{q����BJ�RL��u5�z �{��pH�:��>-~��6�S��������r����W1��a�Q�,�:���I��Zs��4������D���`|\8�b�\"cZ��w`���i��5�ǻF��_SAPgy�7#��	T(W�8 I���ȥW��6�����t��T+!��I��:��#�|Ce0D'�S�1*x��\>���Swn����xGU QIɢ�`$��M���_��ctw:�&(��,e���{J�C=��Q;	����/�� �CCq?P]>�&�E�#������6<n�8\�*���LQ��ߊ���/�|�c��XW���B�%��S�Fl��L����	��;��DFb�Q��a6�����A	��P��Y�� ���m�3rr+.ZF'F$�ts����Ed��)d����.��G�@_�6[V�4�����2��怫?؝�����f�<w������� Bz��_����0�KI���'a��D�<���X�eO}�*�:>D7T<����Ԉ�E䶴ߎ��Нr��_:�_���N���i���{�H)�0��W���v*�]Lk�n$�ϗO�s|T��iR@hx��_�]�(��~�+�:m4-��v�X�	6���tO]�nNL�eoVN��Pu!����䐱�N�X�΍�$��ii����-�����.�m�nOU4;�ɼg�����3�L�E�&��a�}�t� ���z)H�M����;�%6�SyWX�5%�PLv�a��Z�5E�i�{�1t|�M�%�tH�7�i�2����ի���,�w
v@�͉���f~'2G���]�ixP�3a>�v=��e`��9)�h�8�J��T�X�*vu[�˦DUۄ��pM9GT�4�}�o*n�Nw|!���-BT�a�7Y"��jS*d�֝d��#��i��hb2}?Xs���b�t�^������v�ޅP�ٙm��D�z����X�4�_~1�^	j�&wW��/�X �gY�q/��W�F�'F�-�E��+~p�Ϧ~�J���f�Ye0�/��A�j1B�%�LG� ct�)�(�̛�Z�N�n����	�����bģ�l����¶'8�����&�ۅ�Rh�>��,VJ�g-�z:/�/�1����>����J���L+:��~��:��UĆnN�ߧ�;��D��y�����/�0�9U-�@2U_jZ���[|�(#��I�r{�5FqŅ��0!�T�E��R��?|�JR�z�j���|�t'(��\��-ۗ��,�����TIp�g54͕RK�4Q^`W��}n��%�|n�^���,�z�g:��s��]h�TLS]۲Q�^�K�>��V&��+Q+����y�pXw���4�/,}�`���vef���le�d�Sq.6�d�.w��9�G�E�F����?&����&�,ؑD�3�][�6����0�?�R��<r�k8_z>���r����Mf.I�*��!(�����f�PFY{),�tW�{f���w� ��B��䕒�3S�di'?�t�K'*�m��. ��s�*�O ����	�rRSը�{`���:�pf([=����L��>e����g#X���(�[�	�Wx��
+$s����aGN�K>�v�҉�go�9$Nm.?��#�}�a�e��_'5g�� 6���r�p��0~��>ߛg�	�e������:Ae���7�D��*���7R"v����+��7 K�͓e�J���7�\�{?�8+�gW6�&-ur��t�>��{�P���+ThE��l+	�}j`��G�5�s:�e���U [ߺ1R�"���U5��@�]nU{yv9�܇�b`�j
���&h'rtm.ny.J4	l݃nH݋.�/��E����a�\��"g=7U���"���G2�N�YY��=�Oc�U�Ӽ�����I
�/ag	��Z��;�3 K�	�20�t@K�@`+ڻ���?��D_�n�x����b������bí�Mx&���6o��G�^6_���&Vez�-��.�C�Y2 ,�-���v� ��N�Jޭ(zo�^Kۇ�۫
m��#Q~�K:��Z�����:�������"�g?����\�o1�B���_,�S�M�m�K�������3�`�(���L%ܾ��M M}�ԡ,r�'��^�M�]Wk7�ް<%��h�z.P[:�n���a9s���#��L5�UL���Dl��^�F������|���i3wT�X�s��~k��X߮�8R�Hr��9q������,���L�N�ؖ1��ޖ�תp��nsP
�>�Ů�|	`Dֺ�%���n���r�2M*_ ��D��Ԑ@��TMʁ�!�������U�4^$%�Yb%x���~�-�pי���E���.c�VH]���8���P������Ӹ�B�-?<3߿�'���+�����U��Ua��B"RƢ0<R6����8ad��E�g�_&��2��1�05���Rr� ���P��36`5�c��
���:������=R���b��~�pĖ��EDp�p�'�o�J^�ݞ1����h;�? >�#�����^X�����d�.����"���ݸ��BRġ��ܹ�H�^gk�CÆ�hQԺ��M?���-t�e�J� P�|.1�Dq6Gɂ�*�)qc��M�8ո�Zr�ϨM�4��|=�~�z��s�ڌŎ���k ��M���O%�B=TiF�{��d�!$�;�4�_���8��+\fC�[��Fi�͞%���3�C��0nm�%�+�ϙ?�t�����&3��ݼ��|j�+7�c<P#��r�:in���cz&�dw�{����bb����+{e��/ڠ+6"$Ǧy��F�9|=6�̥o,�\]�W�j
N���fZ�>g΃:���\���;,p�-nÝ�&��^���
���U��K��<�S���մ��7eCҪ��d���n''��Ϛ�*��7�jJ\󼺏��;�8��*(T�Ĺ)�e�s�H��e</!�n9�B�P�v�ٱ��đ\�UV;0��9��L�����<�zi4lJַ�L��y>���QhxW7|p�P�k3}���y[D�'$Ⱥ�,����D�M��z�|ґC�ۥr(+8qh+���������N���+�.�RB�����B��=1"�"S����LE��A���>�5�>w�|�%���w�qz�ƪ���&�mg2�⭛F]E��]��	�����4�<M/�!+3k[_^���v��(Ƣt��$�f.v	4�W�1O���q^.�l DU�3��c�f|Nr[{�1���Q���#7��D���(/�V����!��pC�C�.�	M%,fA���!}�"�z���J��R�Zq%D��]��UGKo^TS�2�X�<7aD|$��g5s�CV�SE1����Ʉ*mm��f��k�p�
��;�Ҿ�Sk��,�����v6��ǆ
C��v��������z'�|�)�a{Q�8Pv�M��a����1썂��v���2�pd�Ol���;e`�7�&ٓ�vj�UG\2�%���>,� ���>�O7�VX��c�=��{z��`�����x-�G�:of��}�'�����W�s�ɟy#�2���>	o*���7,J������ܧ�ڂ n�`���]1k-�>��k]���A	T3$E�aj�w� X��0��`ܬF� B�!ZA&�Vid�;�Ai4"w5�2�)K��c���Ǽ3��ޔ�k�1��ֶ�J9,�!l�̰P&�(�2x�f��o���d\��|.�
�/�\�!�"<����i%ݻBiS]ξ�&i�Y�>��X�]䦷��+��`|�Z�q$	���4�oi�nUoDU����7�����y�	��p�a��Q��pܴ�R�n�DI ���
����<޾��j_WX�+Go��xdɈ��uӚ��q���R�
;��yESo��|$ps�Ҥ�7�A������\#��{�*斯ӹ��Eᷤð�
 HC���w,dx�~T�+�}�N�/�1� -Hh��D=p~ K}	��f�&�3j�ó�iX��iF��7y�����j�dT�{*��L�3t��%�a���i� V�L�U�Q>������݈���`��_}���Yd�5��`�#��__M��vfv�Q����Q[U�k��k�^�A�!���I�Q�S�H�w /.J�`5شIc�}�ݏ*�j���2$����W��A��*���^�x�!6ף2uO
ީ_C"Mf�j���P��E�	p|v�-�M�dw��Ռ�9��(��ͪ�]Q/ibd�W6�2�� ��o�������q/�,�(�P]p�D�	�3�9s��ig=yc��c� ؚ�J�&Ei�Fe;O���L��9�G/��R�W$��khغշLwz��gM�����=�p�iѴ���7��J�<Q��Բ��]�(�+�܊Wo�;�<��~�aDI'ݭ�P�J�޷���=h��ϟ:g�y����0r2(�p+57�b���p� �/�H�&���7��Y��j)�yy>��B��yc����U�Lv�Q���ȝg� �!p=(ёg�2�>,�]E���@1�DzI=s z[/`7�{�Ǩ��������
)�2k��c��dؗ�R��m��Ьh*��`6J���`E��ͳ�%M%�6�5u���V�.W)8LxZo�	!��l�;J�8|�QgҞ��2���J[:�{�
�g������v�#��r���QdFX)���- �ܺ��Ǌ���"��߉��Eu��.�kl�ӈV$h��6O��Q%tYg@��˵v�0Ő�Qƭ�Z;�c�^\22��0W�G�fuY��_D�����ɠZ����6Vl=�j���DHu(���y����U����������'��L8������:���Ǭ��8�o��oM�/P��̈���֥b�Ѹeլ�(�qtg����߳��R��ÜX[����dݼ�|
=�0�z��yҼ[����X|U|}5�L��~[3莤Tt�풂D)0��8���6p���<���d�����A(@����q�>56��y��c�P�,��x���x��Ruj���h��U������U��n�|�KԘ$/��č)�^�����d���ա��ǹ�k
�et�nu{�B�`k��;��.�ڈJ���U����*����0\���ut�F��見C��=!��$�!Y~��C#�#�Ӌ�T�*�NOi�ӯ���rj�0Q"F���__(��G�:!�i�u���t)q��}�h�����4�?_dqQ�Z���l�~c ���Su�<lI	 ug�@Fk�`�i_FZ�"wf3�w�� d��p�i�.����	���.��Iϩ��N�����52bǾ�����w̠�*��D��[�.�|�!Ak�S��q��|�Ϟyxw@��I��?�_�0)����y�M#�� {��0�C-�I��"Ŵ��0v��%��zAv}��E�'	aS����h)�-{fE��U���tO@{���hZ��D#�''�&�ր�Z̪V�BWi�\ry�}g�A��]|�Z��r�Ks��8���3/VWIUe�u	���[y<���M�p��ǵ�K[)�r[�h�,�[c�J�`���R��~��K��".� d���D$��*�)X׮Vh������������P��My������~����L��TW!F'�U�����j!�2���_#}���tge��7�7���<%��,㵕9��G��1�i1˼H�8�P��
t�G1j#@h-��|f�U5jB�g'�,n6wߙ'�##�ҰZ�$�*�
�ݽj�ZTцy��i�,Ӈ���ˬ.�ah�� �.q�oN5����!�y���n���t���\�E��g�R-e�.6`Q��|��=�>�q	�&=��\7�k�F�>T���#��.Z�3��߯����{���(���ED<Nu�\ �0��m2͜s'�ŏ����v��g�k���V�V����v�[���O}�`�O�P̊0@_[�ce���
�0!�Y;,�s�A�_'S�����'9��[$(��s+��l@<�m�0)=%�ST䚇�wˮd p��=���m ��(8ßW�d���6_�v��Q��89"=��q��ۼ��9�w���,�5�$�C�)-yN!]׈���4���d�QBB�:(ݑe��z-.�܂�PA`�c��0t��������PJ�>,.��rxTp�`O��5+�af��
'�2jj�����+6$/�)������Tsڡ��Ɯ?r�'�(9][䀷$��BY/�Й�L���[Ġ�{�G���z���Ί�m�t8A�X�+w����\6L�ߨ0�sg
����C��%1-���50�]fv&}΍&�X�����I�V�u��X�n( �\"��Kw���b��إ�v�2�Vs�\��*���!��7o�9#y��Hz�<�[�-r�JM^T�hSʤ�'��ɇ����Gt�̚g�N�47=&�
� �v�%�B�d���B��-3��; ��Bc�Dh��Gb\��+mFzt��틮1e1k�OYr��x3M	FM!"ӵc�e\�(!Ec�&qG�敺3^�MqR�@o]��O��r�\�&��+lK@�I����!9��2rt"������W��1C	v+�+��3(褷O�{��;���VVo��8`,?�*�N�����z�/M+��}i�����I~<�l����u�5��A?-�I�g@�b�uE����q�<ɀ�?�!c��a���;�/Gm��xt3W��oʙ�jvA�)e��ΥB��&N�@�X&g�B�%��FMBy��y��g�@�M��;���q̭�w�-�@Ʉ�P�б �+ �U�"���Ӓ�,�!���ۮ�2�.�����\�?�����"}�"
��+�l�/�V���x���xO	A�����"M��݆�6+���G6�^f�4	�:J�i`��L8�;h�C��Y:�Rէv��L�S~Ќ��Xi�wןD(�,s���m8z1��'�aM���YUE!�ӋӜ��]���48�>��xr��h���$[<��������Y�x�2�B����W�G��}"�;�����;C6��޾��bn�<	�߃j0����E@L}�"�Ƭ.^��2;m���X#v���5G�U'=m\l1�x$��p�	�~Q2t4�'�Q�ٿ��8��������i��Ptg��ю�B�R�'���9�!Z!�Ĉ*u����@4�����q	�Y�j���,�K*F��RPP��M�~�W#��`3��p��$��������;�����{�Z.T�]A�s4`U�C��T7��X�V���D�q!P�vSLA1 r��t��#�J����Zb.�;mtV�x��v\3kN����v1�NH���K���H%�vg�&��ɇc�:�?Œl�Ӊ��r%g�s�9k���;���g��淲�\��50�_��-=o���z�0�����+k!-�E��/*���>�5�@l�ٹ�p��v9���m�?kl-�Z75���e�O����*�DUI�:����X��
�p뮦��~�� ���}{OZ��zwL�[�V�ۊ�3���zn��ؓ{n������rW�$�LͯI��ƅV7T4�7:r�e����X�ƺ��{��%�Fz�T��0A��,_�~[�~8��Ҭk:�r�D�Y�o1f~H��zEw0W�P5܅r8�F;3ؤ}�n+6�԰:]n�/���~���
��U1�@e��R�}ee��{[Q��ϒ���� �p��G�x��Cr��Ćp��P:|f~�I�����K��D��X}GPl�-o��+�`�4)�~��P�M3�sR�\�!s�zn��K�Ĝn��D5�ay� �����s�B+'-d��AN������W��2�"dzx�35�]���%���<���\~n�\�j�|3�!mh�M4����W�鳹�����q׼l<6�z]�t�zѻ�pE&��4���
Y�|�qG�M�/���5��S������D�]_)Ց�0��W]��$�����9:�\|62�(E�����P�{_���4�:]�ngwYH��Dj��vd�b�V@)��� �1�4j�@�w�K���)����t���.��������W4-2w]�&��L۔�6�"0�0��괕���l��=�lɯ�f��{�m�-��:K�E��.�g �� �z��QP/0<�G�	�$�U���y��xӮi$x���^.HeU�ȗԤ�(t@�<h#��*e*ή��I�]�K��V2����x��T��vȐ �il���5�4Ag��;��sHy7_��i����C� 8��	���G�$�X��Gx�u����Co���p�o�a�Y�@!�S���b,���_�Ĝ1בf���v�%L`B�ZP������`V"�F���~m���5�+��<���:,�H��~e�q��ɿ�feR:�NՊ�șP�n�x���
+�O���`�O���n�)�{^:ݼ�ưf&�q��:u*���P 
��
���9,`8#{��͞�{o  M#y_X�~z��.�����Fhg��sKBސ �0����2{��G�D�0������å|�M
3`��a'!RG���c��is*oj��'
���m�~:��O���n 6�*?^��0����V��F����X�y�$O����Jin�p�J}i�����qVn^וɻ����i�<E�+�$��	�j�ae-|���J��I��V�)�T(T-��{�։�xlc���}�I�@�K�H�A�-�z��(x��fy�'m7����eo�����[s��U�0��@d}!0��>��rIa�!)_%�Rvx�˼YHG'���M�P���O4�;�d��pڣ�)�n�;#m�<w���%�)�AT���N�⯨2 l@Bt�君���O��a�S��0Hz,�H�Ig�}N�Rg!�b'Ciu��l�m����p땅��F���%�=-8ό�	�`}������Ypy���<5����J��dޱ�B��3`��XT��	y�|��	�Q쐓�.11�9��-�kÎA����t��ߞ��fB1��������!@�/S�NL`���zڎ�ه��N`d*O���~̎�J���a��e(�3m���F�3Ւ�������&Y1�8�E��`$�d�"�8)G�?Q�D �+p�F;\�� t��Xv��qq�KƎ��O�z�dй0������$s]T����k|�0v����4�qX���|���{u�F���R�w������fVbu�g����n�t[�Lo��n���&�sʘ��$5^\R�;>�~[b��^f�n��'�0�3b�^���0GCfKRys��c�pG�V\��g/xY�W��(��S�i;�s3��⼣�D�|��Ԥ�{��\[te�f1CҎ&��I4��|8���D[�dt�yʊD��;sKL'��vi+�j���zl4�$-�M�2���nM@MD�"_fmp:OH1��\~3ˁ[][3�k�2�AҜτBf���i�Bu"v����-�Yl��̉�@|���>�eؗ�U[�)c�N���_yW�%]�0f,��>-_�H�#����
vJZ� ��F8��RM ,y%�= �7)!�ct�jԤ���6e���շ�f���T�5��}ocT�=��[Q�!�'�D������o�߾�I��	�� ��SI�]��!^)�X���cߧ5�|��x7�Yi 8�-7ǧ._v������C¢͉��zu�h�.�2�k�D����"(E�d�8q˄��`�@Bؒ��M������
}���T$센��8���L�A0������s��`֋Fo�s�}U���6I�^��ʵ"�$�O'�V�1��Q���w������뾾��Ϩ�ߜ���@D�S����Q[���!�9R��0cE���%�W�-�U��>gBZ�a��c�V��nϬ;o�q9�kH$����SQkx|��= 5��M�=}���-���i�-���K�2A�Abk`Ru����V1�%�u&%�ćA/2@C��*lxr����M�@��c�ӊ��|��wm"W�/�TAb�L$Ak+zD��y6�]��5]7���A:�ĩ��{��e� ��|}��Cp�(�^�*J�}�l�0ܱZe������Ś
iz��k�{�m?[�qdcb�ױ�@b((6�9g����?�Xj���ϭ�^����Lh������5p~n����Xd>LD҃��c�M�O�ƌz��E�D�%��w���E)�Vl�.�;�� I�!�Jc(1��P"	�y��������Y�c$Lݬ��E]�t��ؾ<�P,ܥ�	5x��>µ�$&Y����WK����Z�ĵB�뺗�y��?
$-�K����~�v��sX�O3�\qfN��5E;{��vJ.Z���`m�	 r�p�3��".��8\/����[�ҩ�R�J����:0�_'#W���aP6�=`���ᳩ|�뾳����,��Ѽ1��+�D�Ԙ̫�`��2H��c�u�gQ�Ÿ��w��]�82��{�V,��Rݯ���H�p��C�!�g�0��,��Qn5�U8z
�]���v�Vqp�r�S��dDƿ��������y=:�ލ����%���Q�Ƕ�8�`ƙXh��M-�&�7%mk��Ɵäć<�7X��:�P�ؠH~�,�.=�X-������&� �{Z<�4-�
�aҜ���Ĥ/qC�d�
|U��z�5�^�jə���5&Y^}s�7�9�n"�_��I/+��%�eKu�v��&t��3�I�J�
�L$Vɶa1֕�șd�\R^��ߏ�����=�Y�Ma��p�����Z]�1}�P�4��*c%��o�d�kU�Rp2Em��x"�B{�^�[?���n��#H��"�<KM����ԫs�90�+3;��{*W~ɖa���/6$ʫ��$k�y�1��{�p����P���b��K��(X�)E�
���=�52o�2�[L� )�Bϗ+,[&��$��ܩ�"�\AE�"��+4��]�rD'{\��jA���涉�d����@+��t��D�!�EX�?cw[3����
b	�����orr �W�G&��E
LE�[��&�AH�F��Y��k&Kj�/
nq��2ͩL���X�C�lo��2�s��4��Ժ�h��&�E�_�I�:~�xr�;1�cQ�Z�����* �=�MQ)-Z���G��5�̙���OH
ǻ�� �ԋ^���$�O�Y���VP2�xm��	�p�/2�0�o�k�W�>'��������i!b:>�Tp3w���F�l�Pg�S]��~��w�F���4�hY<�5�'��)�Z5�QA�2�L�(DCF 3�!��(��lx�Iz%О�L���4^)�j7��������uR�kwF�d�UOk�p��]i�4�+�m��t�z�ܢ\^��
\��B/D�������p5�"+�\�^�*3>� �&>�?o��b-w�:n���dM�8@I=�����o�����iǊ�LX[�%4�*c�H>��
�5��20�+��暆�]ϸ{^	ٙ}��ܻ=GO�L̐0=���`㟬v�BX(%kb��r�TW�-i����#��D3܎�{< �\��,�t�۰9هQ�BMno��)��<��Y��Zx��LTlח?m�K���&qb>-.r�pf��s��x��^���D)��1�}~�<��j�x,G��-䀕�ŉTK��ɼ��}��h����i���C��e�<�V$�@�s����ȿҘu���y=�ٞV���7�ԁ��ff���I��8o_�=-�3�P֫Q8?;B(��E�.��`������KO=E��q�>�V�<�r�>���睋�[{RTbH���6ph��A�1)d��س���%���Cv�8�E:`2�tp����������>+��L����}kLLG��[E�o)�qT�t�r�;.v�A��$�b/�2WlH���V�.� Y��EE��S�P�S$wVJ1�78�W�,n����Βߜ7o���;6�Ә*1Ϋ��$��G�2c��>�l<���&(�ٙ7�!	��R`ɸ`��|acr��[�׃&��J;�[�$��Z5��>]`�E���腏$'� ����e� K�FC��UM�����7���.x7l�O��M��R�~�"��j[�΁F>v�撪�.㘪���X�%��m�F2��� ��c_�ܭ��X2^&]9Hqy���Y�Wf�vf���4w_[��}ۏ��Bn'ё��0���e�{ɞ��OU�5֛f-��r.O����rU]�l��$V$�1 =!:ؔ�)/��3�m��Yf��ߨ8��ލ�����,��.)��u ���m�h�D'�!~�;m��f�x{P�T{!�@����9��s��<�5�O��h��
D�Z�^^�!�qNp;��A�m��I����=ۜè.߂�Nm7>D<E��E������8�~�u5�9q�qwbf]Q2c@ p�g�������� �4WI�y�#�Y��U#ũNKǃ��[٭���'%��V+//c�Zd�1��%��Ǻ��twJWh`(`�p���v~�Q��`�R�el��D��.
�Dyy����gy(��	�V"3D�ELCv�G��G�/mx��vy�_������`�����1�����\*���՞��n:���G5�X֢�U>�`�i8*[\T���}ك�9�L_M#T�鐅7�cL4�f����L����Pk�Fn�xܴ#U�$���C�����l)u���CXT��p��l�G|T�Ȃ�U��3�9R_ A���X����b��S�OJf���5���́�G�gAᗾUT����5�����
k��Ǒ������~O�N>7C�_�~�/7/pߎ� ��FY/T�ن��L-�G�l�����<u�sv�0���6Х&a�� ���Ҩ�H=Q1�y�|����x�TMG���q�+�Ľ�wcT����M]��y[t���E���Ɠ����=�]���HH4�5��ΎcDo�z	��l���Reo;y����/�*�)e��4�~/[�qk���⌆4'���B���*���ô��8��I�1��߼ ��}��L�(����h���E�\J�v���Y
���i%�� ʕʈ�~��:A8�ޛ��fMu5���F6�H�/�t��l�1mY��2�!H��L'�p:p��)0�J��=���7��7 �����!�����2��LE��Π�M����<�M����g}�Y�'�%��ੁ`��v�s�]�h�D7���o�� �R�e�TסYQ��X~��gD}�tC�zpS{X=(��v��ù�$��Z<w�:"�X�T���Fv��:2�]q��+V�h#]ܥN1F��#C�5-��v`9@[%��z+�NҞ�:m�8[����h���^�K �� d�}�X���Ԧ����Q7j��5ء5nL�,�oU��~�{%����(C����m���j��&��>b%*Ⱦ�XBA+�ov��10�#�����|�Z���D����4b����*4�}�C�;gR���,`�	�o�(�Dٽ�M�\k ��q+,�m����c ��%��b-ڊ;]b���Ls�s�}����UPm�e̲�@��ɡ�s� $�{t�(�82������$�����pT�@���m��TT��q>���l�۪�G��j$�C�M��u��C���q��:�L&k棙�Y0<ܾ��>.���ll|]�� �uY�49O1�hE��b]5��w�B)��U
��zH&q���JhM��'�`�v�V�Y�JjfU҆�|���uꈾzn�g�;R6$j�P�GU׈�?_�<�vҀB�>���J���#�UK�>�x�ٟz^��8��K[)�[�� �A���gM�	|�^��w��x�u�(MC��2, B�Q0Q�n+kap�X�GU��g7)0�-d<u� ;�H�ɢ�Q��L/�USJ��
A�$}�'�2uPy/D��2�$V��+�n�g^�$
��՜����!�ڀX��\`\�c9s��6�����&W�Q� =�{Ss�����P�D��F�~�k�!�MT0�w��2V�dT���ڴ�������XDi$��Rndh�Mat�}Qrf����@g�O�d����
���՛��rŐ�f+�ꐦ�w-��$/2m����_�;6b��q���-&d���f?O���+���f�i�O��EŢ�:�Z���E��=�ɮi勉�Ee�0*BTh������]y<v���zP�LA�X����Mq\�GX=�)�������/�~>xA/��1�.k]����hyE9��r"a��Ȉ���"B��Ғ#H�ba��jMӥ:���~6J#q�|�<K�U_��-���2�`�����p� �G]�ˑ-(i���rDY�M[�u�����Qi�?�*�#jU��yۛ��K/V��[�����q������YlV1`ȓ6L��&�lV�I
7L�Wi���s?9���8z.hw�`
й���-`j�\�کWAY�ř���l9$�d�Nڌ�8U�/�����ͤQ"#T/�
�rr�J6�L���9/8?>�4u������dok��O�~ڰ�����7&��O�]<���W�j&�m6Z��W���KA�ޞ� ��̻4���%dP���ecj�hK��ͽ���� {}ѧ�4G^�Q�����!I���� �_{�>���}S ��f���.�E����ԤϗE��'mװ9*R,������i�8Y�!fW������z��������dЎf�-C�6��������G9���^��h5=�@��f��;1�K��O�LTAaA�\���&Q�P �����p�v��A`�Ǧ���D�� �?1�޷ոO�c���ًv��ݷH�FΝ�p�E]ddX-2g��E��A��` >����o7r1��S�J���a�	gҟ	}dq��D	�GF���ɠ�.;�^}��|�*V�����o�CN.7���\�R��*7`��4ƨ
?�A��V�����C}QN�	�����NX�򶿯�MTl��~�-�m��+d��H�� ��N�׍)�nÂ���N e�������&R���m���t�r3����YZ�e:z*��>9�n���|�_C���n� �3���b�	"�i����b���ͅ�����׺@j� �:k�E�S2�R�3e�}&O|�Em�P��Y��U��V���%��{>;f7�E�o��A���)�G�
z|w��7M�O?�1M�ls���8�i�
��mZ��(�hi���N���������8�+!�& /��4��&b�Ph��*&*����w1t}&=ؚ�V!�J�	��\���UCnj	�m�#Tc��C)�!?At�X�4,<����k�1[��|�P\�f ��dom����aO1^�U8�U����`�5V]m{���*�D����1�Ц�l	͓9�v\!�ѡ�R�1�_#X=q߱�,���g������}2��x���7AӲ
^�P�d|ܫd��1.�f��|��h>6g��� |���[�5	���}L���%�=�_��<��oL�H���j<�25��@)Hk0�g{�ѧH�*5�F�p�[]�2�]T��YvU�  d��"qy[H����t�=b|�ꋼO�}��&�Oіǜ_�Z�k��GAe5@	��>l�d6�ԗ������`H�K_5��W%��5K/���Pm%J(Lܑíxx�x��_,�iZ������s��Q�O�։��D�'�:5�I����*jT+����h[�eu�Ơd���D�O*�ߛ��?�hX�	�DO��e�gf�()��*˳�	����G���x$��E��r.P�����N�PE�.]+�����_��o���{���}S�sXW��L�Ζ^\w��ڄ�sQ�j�#����AD�u\�� �ցD\�ψ����Z�)D'y`�6��0�/����di�t�N$!�	���4�c��Sk��E_�@kEKz�+S	ﱜ�@�x�;��!��Y�F�)�#�&Q��9�����?��)Q���' ��\?ـ�4���B2����sF!�Bp�Cz�����q3	���q�Rz�f�gYE��:��Ms\��:�m07�5X5�����0S�T���*�X(��IJ�󂦝����MR
hȏ�1>ldG�!D��=W`̆��4�@�)�R�b����`<:A�źG���1��G���˫���b��7�����h��oon�i!uN�#��v� "�;E$�hK�C�1��U�����A�Y�*.��1Cא��z�x�A��h�C�N��f�L�{w�Q�ìLF��>�^�<"��L���R��0�b\S��ۭ{����]k�n�[�f<�gy�_����4A	 �0�i]�Ni�4��3d=���CϾ����0�jnl!�o��.� k��ٍJ�_f���BFih�m��Gl�)3���n�4!��H}u��M���.�\Dz.Ȱ���6"@��sVX�er��#͙�.���l��K��3�[��f0J�Y�ܸ����KR�:��@
m�>�v�O����E��n��K���U�I��V����>!G���'��dv�aJS��j�:/�G-�o�wAu�F�����o@��55��y��j�!��/�ayЭ|�v��ۂ�v�ϛb���\Y�Ph\6�[>���ru=�{�����II����C�S��,�RL>JJ�M��Ǒ f{2�}�d��(�W^L�C~�h_�������s�U�I֖�\Wq�o�׏��@�ҽ츼pȻ�ɶ�T�I�z�hC0�Gi|�W����{�Vp.�D����tԺ{�5��9UQ9��u|Q���>��nm�(���e�
e�Nisc�8�іU�����~�. ��h��!�1_�o�q\�t���Ma����K�nq��]�	$^�QR�a{��'UI�=T{ć[(" L��z������b����Q�F�،����Dj�O��B�M�	�(ȒߢRp$;��>/�����zn�#R�@�x�R�#�_�'�("�bWL���;��i�=Sp�p�TzI���|�d6�' �7a��0���&�G�h�d�c$�#�K�d���f���L��v"��Nm���AgP�݄���(��B�g�N��9��fd� 8���5�c��U?J����۲Jw���Y�t9h8:a��O�C�<}EXkX��vh�e�F��[4_x��й.SӣK�E�v�}Ǧ�!��t|��ڥ`�'	�C�f����~ExR�s�4������i/�'�yf�Ҩ���#�I!��җ�Xܭ���?7�E��r7��c�<��eMC:�J��9��
u�"��q�(��ʔ����|7�2P�"��&��-�.k��ly"�֠ph�OHr*��m�<��EHW]���y���PO�MR��o�c�.��K��R����Qa��(���Q�s-1���<����<��Y�?�Jl�^ץ������e�i�E�&��ǳ����x�YZX�q"��+6�9;�ߖR��x�@��5�\�g�A6&Ռ.(�ʦYᙝ%����96�1)�ӎ)����cdd�/(2�OQ2e0+.��͹`e�2�H}���6$@C�R/�?�Y:}��bOZn�Z1�Z��T|V��{���Xõ�.��ט���D�P�׆���p*�Ұ#9fWP�S��(�6c�}�!����c��e�������B�<��|�d�jk�����`���p#��+,mqK��3��i�4d5vu�h�6�>��4Ю��霣��q���Ln{����I~��m62��J�"5�K��u�^����v��s��F�7!5�ZF��� `��&P���b�G�lozy�^@��!R�D��\�ڦ9��#ݹw�>��e�<Rh3��[��5E�ϱW�6;�����:�XJ��
V���4X�LO��Ǚ�8�	���i;J�6n4ibx����Ҩܠ�V��ನ��y��t&)q5���<�E��&C�)[f��ՙ��6u�$�v��+��C5Q�mb�6�ÿZ��-�]�j���r�v�4{��E�h���K=�ɹ��`�o��p��$�1uy�8����=�WM'\��(��y�f>��m+��)���q(�|��bH�R��ElJ����b�e�|OM��~�yx��P{�D���D�#�|�yE_ǐ#�;��$<0����?<����z����N�@����d�������gH�o�;���gHS��Җ)`B�*�&�ޕ�Ԟ5�4��|M�����w�l�܍����6o�I�L�t͗�7b�0�CYy��L�9{���ʤC�i:?���K|4���x�;��mf{0�hL&�ſ��?��_׀J�:%�#���p�U�����J�|	��nU��WJ�F+�U\������	�Λ��*(�ͳ�@���.�iIe#WX�$s��0w�f�-�hާd�������c�"5���Qv.&xؾ���\�#)�g��5�Ϡ�`�9=����2j�^u�{_������Nes|^��߁|�����*X��8Lg���Ws�+q�^��3B���%�
!��@)E�[�;ԬT��5�r�m F�8H9��x�0�a���uKG�����*�l*��r�B����&�^��_�s���X3��@/kK�Q�?����W�X>f�I��Sz_~�CxV'{;=�����Z�r��4?��ur����3k7}�J~��jʋ�✪4�kejH=�a����~�3�d�6<>D�j��[󇳸>�hI���?��T��B����Z��<�L�l��'?;!g#ݯNZ�T����؝2�B\΄��ӯ��o,�ߺ�ǃ)��r����������Ȟn߷�����c�{.A^����7�v�R{4���{�����'dSɣS�~�7ݎ���UŘ#�:bX�	��f}C-��ڮ�5�T��tx����.O���j�F*�\���b]ix�n,Ͳ�鮉'��Џ���A��� �PK�t��������?�����I~kj3
0T&�RuI��i)_�z�������<�DPw򂴰2���_�[+a� �i��o�5*����Zlʰ�!��an�ʑ ��/�.��6�BkbE}W�V�Y����^uq�Ewr�51�C��%n��H:E�S�������\�j�}�\g�vz����)�3��Ϧ����T�L��{=�n,F�q��v�l>c��;FҞPB:���2��A^g.'�m#L=���ޑ�ձ�Rػ�5��	���_��F�N/`��)���ͿY����)�=Mp^��=�
����%�+��B�^�㪥��ކ�9K�S��/�"�5�
�I��Cs�~�+L�;��q�g�T�YR�Tj�%�#��Y�����$I�#	�6?�;������`3.�F�SU2�ME����t�iym��\}
��N��:���T7�e���lv)�G�8�3�ʏ��L��X����~���ŭk�q�Z�N���<E��/�䃢�A"9�ű�A�	���Ĕq����YI��PeU��Q㸕Az��aݔ��Z
���l�$לa}�%�Ԥ��H�����k/���,s���1�fZ.�Ճ(%��\�qF,=H�ϰ)L�����p#��7��@!�����S�������������4�{�d�����{n����b�+Mxk�p.�s����-��#;h��N�$<.� d��g�s9�@�8[�3!ŏ���-��{G=p@N�c2��$ļ��2��io�hС�>�H9��]=�r)f��h-{�I��`^���vX�Q�����uyw8.����?�/�����u`�n�kG|G�*d����j!���ՍE���=ݪW����
�ߥz��O�cǘ�e:[I�M�]<n�Y��D��]g�>�3F7��;��6<�����Y��p�K�:��+�4Ye>�a��T�4��Te�BX��f\���Yl�L��v F)r^��H(�G�!����ʬ�*#���@�ɘ �&���>?�(��\���P�$�H!2��P,<�m��b�h��j�ؖ��P��>LS�!�v�%�I'����k�3�ܡb�}�,p�R2����d�R�4&�yT�Ē$���agV[l��I�>[�ǹ#:HU|b�u ���ɒ&RE+��V�H�D�TM��}�	RvR��^~�ܝ%J��ߝ�̏̂����g�}��8=�bnk� �:qÇ�YP;mL�ŗ�\շ���	4�i�#+�WE��
��gE{4��z����p� ���&b����=�����<n����e˃�m�P���&���D�+Bj�r��i����{&�lѩՐ�;gq̋Y�Y{8��<܀ii��2��8�El�B�_qDG���fS�A���X}��Ϩ�2������
�8��s�U���_ǥ�<9N#O]��ɐK]�)^�R�;�>�h�C�1y����,hg6E0c���<5
���b_?w�n�{6�O�:�,Dkp2,�s� 1R���D�
�L�����D�{V2��<b=��Ƀ@N%g����?p�}`P�:eMIf�^���?�5����6�}̮���t\�񍾸��\҉�ش��'���)z)�)���q��T�M��ئ�����{�W��[b��&������k�ҵ���`Ϫ_İu}{�Ϗ���ݹ�Kd�v0�����(�ͦ����z-���?�j߈����G��n��/O-�'妥l�;�'�0�T�Fc�����+��؜R
N1]��)]R#:��m�|�����E�Н߻�)���2�|�H3l���"��L/���fF�N�CTTE�U�:j@M?EбD��9PB��]���?�0U�Y��Jm9��X;��7h�&�� �R-�u�5?�����7��Z}�o��0q�l�1
� dyy�3H�������M� ����(�1�t���I`)�U�h[YP$Ph#䮾�����_��.��j84�X뉔e���g�!�/a���u���]��3�_�h��X�@��a�[���Myɼ>{q��}�,3��$�^�wJx�fBhē^��~�,���!�T���GK4��[����P#����yg��Iލ�־ֵ�^������#��<,Ͱ��>?���������\Swp�\��3�\���2d�&�=q�F�a;�U�)�*uw��/T�]�ѐ?Ichb���f\������5K�q,�+�l1����j��u'/�������еa$��/�ɞ�D�v��Ɓ���M�`>e=P!�h}��r$����f�t�'�~��Q����R���u�?5�B��4�;ꂫ����Bv�Ɩ����(m�w.�Q`��W+�Z��b�Ģ�HDOSP�
vV�9���S9�#��j9�mdÑ�i�?|��t�Q���`�.�_�)Ἒc_iLV��_XΥ'�g]W��*��0����ү=�0n��/�v�lf0�'<�Td��]9%7�I4��/���	s����lQh)�|�W��- �k��}e��M�7�����]^a�`���/S/�·d|�o~Z3K䒴�Й��p���KށU��X(�x��k�4m�h-�YZ<�^�bP�hwG��������֓^BnSS�٤�O�4G���r<�6�GNԓ�B���RZbKC�>����� ��gF�b���&œ���7h!�2*u>�#�S�#lM#�����,�"�_���Y�3X1zx�t�涥�T]'�Q0��[�R�c+K.���E�BI��ŏf)�^��p5)�&� �8��E�FP@ȯ4
3PUQQ�%q��9�bUXC(�K%G�+�e�y�VQ�{O������p��C�w,�����K�؛{���[�h'F>3
2#����$�N4X^�(�o��� v�����d���'_*8�n�� ��}�}A%���=�@��<�N"��=e�*m�k6s�G=N��0�,��
c�lJ�����3v�)M:׶%��`���,�a��N]7����_Yq��iR�y/"��'-�$�s�[��p����LPCA_�m�ӧ�6j�+;G� ��3��m��x<���s�#��s� �S�h~۴m5�������������^���t�Ѱ�ϖ�S/F���`<�`F�T��ǂ�!f�%��i#���8�>]�z<Xs�H��}k(���h���B$zn�r�� ����URٺX-Q7ۖ#�p�'@�T�R]�sM�cP^��-\
�EH��3c�A�01���MO��%co�7��Wj�蓭s�غ�`�ĸU]!A�*1�>�Z�4^�j�X�4lǡ� �t�{d�=h) {���!z���rN��$<�r`J�7V��0�B�<VYȨ�����W�$>p���p�!��&�5L3��
�-��D�]�6�!$��6����y��[�1V��̚�ԡ.nb�t"�(�1L�⮟���I�ǻ�ZUH�m(�i/�����AVGթ��10�X���c\��_t�+_U �0��Y����z�'-��RA��I۰��[�����e�j���
]�b�/�ǁ��i���%��*^���v��Z����Kg��J�ڠ
�
�(�0f�,��u�&���	{E/gǃ*0�|_����x� �.�[�<W�8\%�:��䋆TH2�^ޚ���S�`�v,�eY�΋��f��b�J��\LfHºuX����ܘ��Ro��M�=oP;�L�'b9��	� ��5�� �&�f������<@%u��o�?�k�!�P�w;�Y݅��W�*��aH;����WQ5��	��[3����ZvMi��>k�� �T���d���>����}�#�YYX��=LӸ~�1	!(�E���C0�7ap���S�A�'4���,%,�o�u<���=vr�� =s��ࣄ�B�Y��i�͕'�r�
��F�O�A$A+�1�;��{�Ӳ#>ր�![�|t�柺�!s�^<AWsO���%� ��y[r�f>l�H�쮍=g:i"��j5�b7$�f�= 
�"�a��6e�a���c��;��)cj5�����
�_M<�k!,d��̪��>��~1�
�"*��e"��)�~a�¬δ�ǧ���#�5���ص���~L{y}��rwC&
5P��C���6��)G�����+�J�dw��;�k~'��]T�-K��+���P��Y��H���YWFLNѭ��Fع�x� �E��ue��B@�mJ��q��D�!ˊ&#��XVl��1���'��d��u �zJȺ����I��C�]M��zS�Z����n����q[���[�Ҳ��� �c'�|}���؈���ϭ���`l�R	��B��Oso�u��B����'�=3�A�t���"PW�6i���gh�
Z�æDb���ծX�Ġ��|�{�d��e�S��r�cb8�Du������c����)O�'+~�58t�m�(��p,��d34�T��(����k��u���fW�Y̾����T�y�׺D),^�z?K��[��Ic�6�N��juj~#o��*��@`_�g��Zl~�U-��M��&&q��I�xe�JG��}�:��1�K��ڸ�:4¶<����A����7�& �i貙ٹR��@%�y�˲���z���XӋ��i[���	+�������g�����p������Ĺ�9�0���t<��s`@aa������7�
�85���6C��娩}���%/�wǶ�t����J߽U���6�2LkÍ�g®��~�w�rp��}�#��?�p������k ��bgP�y;/��@hKbp��&�~�� 9�[�aq.D)���IwW�I}� �ކG����{A�t�8�oLC���6WYQ�����*D��U9*|��F$)���&��L����Q��A�m�G��:�=�s��8�����U�߇�4^т���.��j�ʇ���!��Ð~�Jg�����Svsf�b���^�=l2Е}���#����]V/Ȍ��Srz	_?�O��y{���p��G�����崟͝"�ͯ4����T������A<d�]�����f�7�٫m]��$1��5Ϙݞb�Ι�{\����̦�mށ�ŜjC�Z}E;Bڊc���y0�D+`태Ѷ��:#�e�����5J� 'K����IqpU
W������M%`��r+��Q��k1Ap�������T/)��{َF��+���&b�.�	�7t}�N���!�ӟ�d"*q��\�u|A�����Μ�PX���-�7ϢeţN��ɪ�y2s�yŎ;� 'CfF����OD���b����d����d���[�W���?.T�o�υZ2:o�b���CS��P���2�R�Z�.pu�P�tr�ŕ� �5*63�z��'�B�vE��SL��z[��Q�ǘ��ct{�	lI�|y��$���!ۚT�m�˅�x�{Hqyׁ��ā��q�@>C0ҚM͐ٲI��V)���po���U��"���o�0iiQ,��Xg�Z#I|�4��[�|�FU�W�I~��$�6���B���l�-�E6"�y�_�B�3-hs�r�*�ًU]&�jQ���ķo3��> Y\��؎)��$�+!��!�����ȸ��
����B�oʗ�H�	��G�n�b؟8|G\XA^�`8�i(��:���G�1�"D�d��Zk,Yu"'�E�T�z�����I��M+��Q}�'�u�joǢ��v 큣��g7Ќ�����elRKji����Mጺ������z&�b�kZF45�'(�� ��}�ɰ,��x�D���!pԅ��tyh��-Ka"�u��ϔ��ˬ���n�_z�㐯{�T���=�� �g�X�80F�N�� ����w1Ȩ��Z�2�����9��d�*9c(q�/�j��d�	fjkc�O�����5ކ!Я��\�8x&C��õ�^o�Sȍ~SH�;*x������R�u�`*�![����iJ��M4+��1�,�u���p=g ����
�� *!����9���Z'|9�=U0z9��Ta����U�mc�a,�'<�K�x���_����yykd� 
(�zn��9#��hI��)C�c����j��T>������}"s_�:��[��M
}�Z\,b��ԣҧ�񶳵�3I'��໢�n-���7+�!y᜔��B�C���(J*ĉ�t��� ��Gv���x�X�4�e}��P�¿(�O����ޝ��A�=��Lvwaz�`x��i���0�z�@��录M�`
1C���uZm�\"v��M�,�6R����sK����l��Msh���Iţ�h6��e�g%tG�TްU�������X7��l�(rZ����
?�R�9zL�-�5�&��őD3I3O"ruG�`ovS?إA�p���a�ɨ�?z=���=[""�^���8ˢr�cY|��V�X�w�	:TԮ��k3ұ�A}s0�A�a�ÓpL2����6;�Tت&=�;8��4r���ZU��ယs�U�N�#wd�16[�`߄ڏ��h�K�֐{=����_�ǥ�߽�T:XKO�}	e5_���6��!�b�!yX(�&׺�/a?���JRr$�:gËJ��1}�e��$�@L1��g�	�f������Å�>�3��a#���6�)`�d�ϸMK5��b6���fa!�̭+�4�x�]g��S-��-�f�W���zdM���e��6�1fه�v���]� s�x���.�Ǩ�sTf�
i�t��8��@�6�j�b��� �7[�H��/�{���%j�\�X@�-��8��ۻ�5�Z9-���8J�@�5{c~\Լ��KĂ�k�(6$�}����b(/a/��r���眏?
�N��vm�]B����B���к_e��	%��o���혋m��Ȳd$�����=�����?��w}
^`Ѭ�5pV
��x�+�kT�hil�ۣ�AoF��qX�6	��p+�!�̡���u�,��ɖr�^��TQ��_���(-+I���Q��@�3:�`ɬ�S"7?'�<������E�g��l�@���0���w".<�+�b6��55R�tF�_�W���Y4=�G[���3�-�����������Z�S����t�{\�FG��͖�T>Ś���ޝC;�'�5�~Wő�fP|Pi��RL����r"��)~ei߹���ĶM����4=/���ŧ��O�����`.�ak����!�&�yPfB�m�K.�I����P�f�vA<aI�r��XoS��ER���FV9Q�5�,�H��횋�;�όX�s�	�gg��hLO}徿�#k}����)J���3k����r%Z|������9%����d�nܩd�\���N�'���(�;�0���m��>��7W����]v�{����o;��G >�\B!�{(�@c�&�wQ�{�]}���V{Ywjd'?-$?�� �^�����5ܛ�����H�}k������j��q�#�ޯR@��y�2�D7�y�%�΂4���9�m�:ʊe��Ћ3΂њv��6��S?�D����{�M�7Z������:�&+��O=-�!���ďiX�~��F�g�HP�E��v�l
���v5����-�0�Y�5e��tX�J]��֖�a�(L�m��A�0qᣠ �,�K ք���S��R��?��'d��U!U�1�CR��"i�x{aBt(�[���
�?W��,��m�h��R��;�ܖˡ��|�1���s &X>�"B���~q*���O��Z���t��� ���'�{�aO�����A�]X�xr���T	�����Z"!U�ye�@�o�m���^O�FJK�Hv��!at�+^��׌��M+��g.�ށ�7��H;{X�ۮ�J$n^�f$�H��u,�a��'�&N���wܡ��c�A(��<�dٶ�І8Kl$�d�x��$�PH�	��,�d�~)m���y3ZS8|�c���C�}p��c |f�sS}]��`�WǦ�o	F]1��&~�	� � �.��r�o�,��d[�����V)�5�܌s��|QP��6X��5����m�X�P{��Vx�Q(o\����y�vi�ֆ�Xu�^G^g6������
/Rz��H�p��D�B�Mr,���0����#&M�L�j��Ѕ��+�I��Aڨ޶��]ر�;���~q�"J*�6�#��|�%��LӐ��EMݬdAK�\��U�@OR
's���*�+��Z����@;��c�9��(�f�:�;���k����.���c@�/�q���̩)5�3|<�C�-(����ފ�o�&zgg���[�����>9�&�pF�kU�ne�?�vҏ��G�!Z�^��fP�SiГ�C�Km�O�xb�����g�2�G��i1 �GQ���,���B��m�#���xPC������sp�O3Re���R���Uٽ.E1����"�^6Y�]"̠q���Ys�B�&?�ë�2��T<2�ý.=���È���γ��L`� I�c�-�2�ޠ�RIw#1Y�b�ë|e�	�k�b��"�ۡ���,�:�]������g(��H�8���*)iAz�;o/��˙��(��'�V���)���=�=�&����N���D�	^�b�A�ey�|�[�C����#��SC�S�����I�����K�
�����?�9)�]��\��1�UN�HeNxv���S���ݣav'��~ǫ��~�j��B���7�dv�H2�M��"mY�v��:����P~�b$�j�J�nd�V�)��@��s(}0�*�{�UnN@>�<������
�"�b�^7u�{�(�SN���rC�\�̒{B/���ǐFω�*��2�٬�^�S�s����`��O�[��؝Iz��t��
,�4������f�QD�r�P  ra�M���i)J^��Gl�A�S�EA:��>��9P�#,��^5��D+��e[3��[}gR3m�|Ir�$�F*�2�Q@��c1��R`�3`�<'��BV�/j6p4�ʝ���\5g"�_sV��f�e��YZ�lD!#j�A��M>f����V�¿���{��� 6�J�J�V7B2��^o�k�gձa*�%m��h���=o7��#��"�S4��l��F�(�2,�CW�z��D\Ε�>S�Ȩٍ��B���=�6IٗOG�rD2��{�<1���+�g+t��*�%���HqL��|8d�0Z�ѩ�����p�*���☡��Ă��И�
 �_����ԏ+ً̊�����m�dSN@N���ĖЉ}c4"�ǔT(4w��B�|g��Y��C0�_�0�fLܐ0���OO!Ma^��G�'MF@5���$��
�mNk=�C�%��"��{  ���4���wR��Nױ_���|��n�*H}�`*�h�3�u�2��
������l��@� Jm&��W��N*d-�v�Ľ|FՍ?������������.L\����wFj�ؤ̀�R�ְB��֜d����kђ��5�N���� �l�P�Z�
M�+]���� y��_ T|�����h�9���\4�T��*�9�nV6W��@60qb;n���~dٌ���i��_��L�sR��W��a����k/@�x.H�̩�,�P/�K�\�� �i���J�*>#�A��M&8 �7��@���'�E��E[�XJj�-���i�ok>1����NR�V�aw蒬�7�Q-h�c��:9�.	�k�h�1���,��i\ f'��<��b��	�8�|���3� a��]uӗmP`�$���S\?�2����q@Mn�P�������)�����B�C�p���85��|X�x��{�I��]��ʤ�kL0 ����0v̬�~ܾ�.��|ZXځ�d�貓0�/���;�%�ݝ��w_7%|�:��5{�E��^G����ι�͑ܥ ����zYp�B/m._�,B6
�/$F=h�^���ؐ���CQ$���'E�/o	�f�x��إ�!֟F�*Np-X�Z���PRIhQ�їF�/�!A)*�
���5p�v�N!��(-
��\�w�AJ�)�&L��	�.0M����Uvr�`�LC�� �1���R��h��R=���F�R�Q�\�u1���uH�a3&�-�W�:m;����Pw���7%q���Ĭ����e �}���g�MEPb�v���3x����Q�m���_�em躽lѢB��H?*~g=����V�PiG[hX��l=�gq��z�`��q�N�+_=Flq����@0������gNK�L���汃f�e�*�ʅpR�7F�K��T� �I(�0ɧDv��}�$0;�p>knI�b���ZJmH��0uN�KQk��ܕ?�_P:�P�Y�E��h�9]r��o��7b�&��m 9еx�N\E$�\I�vpN�~�l:.;����Ga��K"�<��)Ӆ���K�f�9y��ue��hƒ���{�f��G��Fq�ѧ�Q!�`��#m��-����j���t޺ݸ��_��a�I!m�0��xJDeN��?��lS-����������2����e����&+�s�R��$¨���ڏ�B`��}|�V'G�7���+��}�,�s�}w����E��F:�����JDB=�LR>)$E���) ~�o����Q�tة,uŭP��K`�T�I۪,/5�i�K�>S�XvK����:��֣N���R����0\���^�cqmRr�C"�AI:R����PWv�����.\[������Ә��%�@4&S� �I��ro�X]FXiX� �׿ا=x�C�u��k�ͩ���1'Kd�v�h�I0
�b][+����Fi'[:�����yKѿ`��'�)�%_���{NV�4�Q��]>�<=e�Z|�vo/'x���J�J�\�0��yl G;��e.��)�����eµ���&C�p��T-�u�Ѥ�"o�p���9�\�@��u�i�x���s�;bϸpS'� �[0����ٞr��i����9���O��Т�r]"^���W5nH2�Cko�3���Z���]%;Gl|���+���P�W��Y� �p���7�޺=�&�k��Z��&#���le�l�Y���.��& 3�R��U[���%Z��j�'���aa͘8��PD�
ďA<���͉��߻�;4:륊C���θ�z+����|C�Ԛ�.�Ђ��ٸ?n�dp\SNU��x�JA�>K$���U(I��@Y��e��#����j"?<08���ȌlQx�!�y�vc�D'����1n�&���+�!�s�Z�_�eZ�옾]i��Cw�"v�R��}�'U��<�~P��9Z��u��mZ�9ȋ�~O���X
�j��ϕW�Z��0�:�Wes��kg�9�!Ċ�R$��H�P9�I�lA�s~r]�	��E*��=m���@��(���sY3p) '8�\�}���yF����";�PlT182F�瘋
�쮡wΔR�}2��+��EP����@����=��$���z�۽�c}�Q�N�}7����x�?9��=
�f>�,�+W�y�*�n#�����,K��_�����e��L0��\������(y�U}[t�F~���2eғ�Ջ���Qa���r��,���u���4Qĳ��ǻ�59��'��ɐZ.��M� ���d�<�y����J����\*�������Z��_DsK����l*�"/󬲕;X�9t��Z��o�{�G��	���Ƨ�Aﭛ�#��Պ��^I z7C�J!�HK�Pt����y�h�-˻7���a�_yKT^9%{s���Yu.V�oA�%Нmt2�@DV�YA�;}߰ؼ1�k�����j@ӗ���^KJ� )�V���e���L�1OG[|Ң��{����ջ���k����\%1\%Z�@�Y"N%ɓ!�Y�͝�=O&���q�LV_N���?,8.
�ECZ������(��3w��&��~Bn���~	���yr�]U_S��5 a�/cpb���Z��q6����W���wح�`ug�h�D�dT��*�����]�z���r�D�^Ō�G���]���"�zn�x|�%�4��q�/�����k8k��],�����W��Z?o��"E*^��YD�\Y���8��c�ĉV�4�[�`J�rI�E�f��a����M+�����?��VН��z�X}��y^�&���yf�3�/D�}*�h�������6����FS�r����>��� m��VBT��^�٥ߓ���Hp4�e�Z������>U�ϛ������L�n2�m�v��~	P=��%J��6�Q���0l#@�&��֭E#���L�h�)��zar�`n;v�Ĭe>W�* ��X�kZ��f�te�T��j\v�|����\�=���D�9�hT�-8�Sv��@*�����ɉ��Z��c	��[͸��-�@���Py�$�!���2"�Թ%��eN�K�_k�O��S���i��W��?�`,>0��1��^y����4M[�p� �@�4��cvV�5�q�H����IN}�ye�T_���W�2���0�Lv��qR_7q�SQ�$�p]S��Ƹ��f�%.U����8�=U������d*��4F��v�+�'t�r��B�����f�J%cɃ��$~n���x(;B��֒�.@�,B���*��
�N?�r�Xd��M`�}d��#h5�O���W�~��h�gH��,Оd��\u�1�A�`۫9s�Ma8\Vd���/�~�R�E��9T���y*�9ٗ�:[4|>����ʂ��.���&ujM�����D���K��qj�\�Ի��n�\�r��G�-��H��������E�juf��BDہ��'u�Y���(vQ�A'�qA��M�h�؟~�nGb��0��l|a��ހ\.}e˒�ޙH_��ztH�fK&� Ʉ{ʵ�I?�n4p���@N����=��A����{!�o���B������E/?�g�z�XJ�l�Oѣ `�K�����<\���%�eC�u;8��7��a�ө\;C��?��h��gީ*��C+���lSov�" >�h���S�݈�k�|C�OQ��������7����Bq�L��D�^�~���t*��Է�1[x��j�*�����(��18ȅ
 �����,w?f�c_���I�(y��[��s� [�}�h�8�u�Ծ]ݤB���pX٧�fb�:^���U������5i ��J�5�aQ_nR���<��n��&��l���?O���\���c�T���ą��n����[�.��}Q{��7��TND�I� �>ۋq�C���)���X�9���^	��*U�p��t<J^�a:��o��ґ���An��3�Bo󞶕����O���)2��oࢴ������?wؙ��Nh�l�K��CwAr��{_���W�l�I&(�ʶ�L��J�Ϡ_&�GD�Zа�t�8��$�Q,W����W�+o.~�!��R����������$����D�1ı���<u%�H�Ô�����o��-���t������P�x�A荋7V/Ps��	ݚ1�p�)����c,���U�0|@Ǚ=��r�h���գ�wt� �[��R�	�=��(W
����S�i��>wP��NrW�o��S^�����I�GA���H10�ǩl9b7 �@2�Z	.`�Uh��ǌ�~R�6)F�0�	�V�TG#-x0~7�
�K��֗b����:�>
�N8�
�7�0Р���9�3���@h��ym�ti��������u 9$��9�kGg(�6�>���zZ�S��_hdP��#�k褝�4��L�N�g���f�E������x_Fp�a^[ߖ��ϐ\�KV�*He@H��M�����Y�*�08Q�	�1⋤l������/�Ut�*T�Ϫ�ճ��ؓV����8�a}q'���Ao��R���嫔FH��#�%t��$#K>�2s��@i�_�ݡq��07 rav��r�G������_�[Bo�#��Y�Q(���)_���0�)y嶋c���nѦ��R�PޟB�_p��Mϕ����*�wJ[�&I7;�W�rƔ� o0I���_���ĳ�P�a��"�Y$��nx&Y�Kp���#*�ǭ�!��S���`��->��UMz��86lχm�%_K@�DM` p YR�Uxeax�$2����ӧvB�RS<T�6�ܚ�#j�:��'��Y��0Հo`؜q�8;LN�?I�� �?�WD���z�+p[I<�}���ONs�'�>mѸz�X�h�/t���0
u��E�|D\C��,#�-ΐz,�V1��;����m�3�EV��C�n}����:M
��z;�9WTc�)U�+~E�Bg0Q���xEƵ�O���9�7q���!gk��3ڿ��c?j �<l�Q-���o�$f�2���Å��b�Ja�=Z��uu��ZNz��H�3
��H�%��k�����`7N��0������x�A�pTLRK��(F�}��A[�����"6����>���6	��ɗ�1X���%�Q�w�YT6��-�4T
��6Uċ�;��}5�L�`o��8$�&T��+����Z�S��x-���������]y�w��e����(��r"1R��*�����-e?�.�u��
��&TPX�\��l��+Je���o��|�f-��,�B��E�ŏ����uW��?!��%i�O�������:=$1ﭲ����K֟DG�$h3J��
U�)o��zW�\3�1/4<���-�������qi���t]4"��D���Aw���v�,��&�ػΓV����ۈdCa���۞"�m_�H�?�Z�|RY�/��*�g
|��DP����==N�aq�/f�Q�Sa���DvP���xPW��S�E�G��W�m)}�4lY�d��sk�eh:�x��'��Vv����e��
��#h�B6|�>�y�:7A�ق�꘶b_�)`q��c_�߆N��Q���� uWQe�i��w7�&K������U��"�Q+mB��am{(�]��T$X��Uo�i4�x����	�^f��ݘFꅭEZ��h*�z�r���b3T&N6�z�E�xy3�*I���9rr�C<��koR<Y�w%hvb�k�S2�uy�v�sW��7u~��a<���S�̴b0��P7���
CX�ll�R�Ř_���H^�YflI�����Ұ��K�$��v�$�O#��q�h���G�ˉ�@z���o�E����#F~H`��>d�^�-�鑼�Wd���:QAi=���ʫ/
8E~d�!�U��.@�5����V�̅*(tV3R!���F�T�O7/���z�ĘG}�i_��4'T9x������Y����*�'ϭ`Ј��ƚC�K�z��T���i��^9��ʺ�V2��E��
� @����n8��U����愶]D�4�D�5a�y�$p��x�f�/�w0<�-�9�##C�z�QWFM�Lc�:���R?A���N�NΌ����������7���W�)a�ک7�k*G���t�5���]�Zک�Z1W���_�W�{��h�[�cfc�i�Q
H�a�FدW�j�o�:��1ІE�����u���ҪP�#�y��4=��h�����&�!_�=ޅ�ւ����|c_o�q�{�h�z�����h�ve�3cG�i`�㽲؅y-�����U08���;L:{*���_{Mܹ��z��0�Ɠ=��O"�3B�a���͝"��y%~3�`�ީ�M����8zO�!�W�g��e_.j�h��$���33NY^91RW�:^�[%M4Y8�^ðS҈�:�_C_{l!��>�`\�,VhͬH�����¼0�}��E�sK��@��3��]ZW�*o�3�~�:D�:)e����K�x±pg \b@58��*o�k��%9����Z\���|�����o����#�,Y�2�<Q��#�p��qj���D���FOA8M�ׯ�>�y�� yt���m��R� ͑j��a�� Ǻ�C��s+]Q�O��!V�}��8�[��͍�`Ո��Ք�v�)�`�KY����~��f8|�U=M;��{�q7e���g�����A*�ov�Q��T�`d�>/�<٫��� _���sx�����":R���+������'a����
��X�b� =��޹א�k|�Ns���ː�P����v�ҕ��ȹ!��>�f��G�X�#���\u�	�{��7�N�\�H"�o<��P�\8��y{O��c� ���iX��/�mE�^����9��nv:ֻǊ7�Q�5�XV����T1ޏ�JG����xp�ŧ�z�yx�y	�1�eL론k�xU@��ãX���F���w���h�Fl9�5��;��Y����n[C_�HMifgĺ�?E5����<�C>*���4���^t��L+�'J����K몳�t��ߜI6}���҃���Xp2��Igi�v���`|4ȴ��ҷs�A�P����--M>Txx�|jheA��7#\�qK.(,�c!���m������:̫����(����ܶ��(��Xu�KacR�Mo�>G��K�he!��O�^�Y4�D6&����_��;��FPU�q�%ob�	�̥#�&S�,Z�ù���lڙ�xP$��L�ő;ߌk�Zv��-u�J���w ���ǋ�TW�O�*�Z7�al�W�/��,>�G��H�^=Ѹ0tܘ����O��+q��V>�QM��mt�h������f`���j�E����0�%?���qbƬrC1�6�(�姩k���ċ5|D�7�pC}��}������ز 6����m����-�1N��#��ώձ�YF�9�7��e��+�E�5�j A���S=�$l�����]��P�c�	Bg���4�f+�����pm�/G�!��b�
���ܹ��Ne����$�E(
K��$LK�n�su�:ȵ���T˜S��Y}n����
U�0�8�>J�x_&�s�������!�O��,Խ��[��o�UI��I�¡��X�rF��d�!�t�%P /vN]�� õ�wIJ�
�j���"�q�y����_��~`�0�3c,�=�mT曎)��+ "Ά��2�8J���[V�hd �.�qS�?�=Ǳ���ck)���N�6.Z%����l%��}��VX�=�%���:号i��P���Y0��T���� u޲4��ǩQ�ԲYl�Q��}��X1�sǒ��λ-Ә�CZ/���1@�l�uբ�&$/��X��{�X�L���\�ht���� ������=-琴Z%&�4`+���&���H�3�Xi
 ��FE0�Nv�ٕ�E;�����? 6�<>��<�?�ٌ���9����a�	�����n��,�sLЮr����%`�&��%����IH�+���Q��A�ab8�S"y�ݭ�Z3m���B�n ��F��W��x$�0��wM��4ә�#���7Mu����1Dԭ��Itu�X-���Hr{����LKAqƸȇC�sm5-(���z�::���]��D-"����3V���C����q�����?=#z��B�
��Rd��N%�
��>�\ 阘M,fo
�ޱ́�����,�?�Gl4�f�>�+�v��^[�ا��)n��An�}�mܮ���8 ��)?c�0��]���w³%�Nӓ0���|��x�܇�n|J��#^���H�J�����7��Vߺ�U!������$�oơ��k%�k[;�@pw���W)�ȫ�^B�u\��%1Q2��یWO�X��>8<����jW�L�?�Ҧ�9���uۯ陘x��i쪬ׄE���'4Z����$Y,.:��v�?2hkn i&�<������
����.���I�DᲗo	��K�kVd�3� EY�A�e�,��{X��D���k3m�]���RQhĄ��r9^��U������)��-kq�zup�_e;�	�&&���;6n�x߄uq2m����������<`� � 8��kC<.�^ �C�^�`#5�3��}�^�0X��#2k^��ܻ�y��s�z��̎fy�F&H_��uO�H0JG[�|����&��P'�^	j�- ��]�&���{ �h��«j;S�9��TFk�k��U�N�p�M_�$�iw�?�� �5(��{�۬~\O�V'[���+*�uρ�����i����:��a9鴛����ƀ����k�2 Ubp㹩�վ۳���	��Ɓ�UU�4^kkT�)�sr�=W=�O��`4������S&
��O���;� ��5�i(�>�v�PN2��ۊ* �qzX����.``�1	½���/L�z�{�����2�D����r��i����ݣN�[%{%��h{�J�gn`VI8RQ�N��#Y��{�yM)r(��k�~�q 0rKT���ud���p���Vm�,.���6S�h]\Qh�����G�UvZB�9�.�(N��ظ�)K:���g�-���9�_S��;}
�oRG�3�Q7%��	2����^�����g�́��5���G�e3t��i����-"�&1w{�q�\L`�����E�V��Hvǟ}�+��L'_��i��|.B4Fh�A�?1���a��:)7�w��g_8"���@u\�s)����%&zw��pa���
W�$�jpMә�7ǌ>�B����1�^�R~�&/��V���W�<�n�m^}�nx�:��{�4�J���9< ؚ"ȏ��V�J�f���%?P_�)BW����0�'O_y>
:�d��1 �c��$���\#���|Xǹ2Y���2���z���Ⱦs�J[�c]=�:T*�
�:xU�&��%�7O�[�����\~�X��1\�G� �(T*r��
�F���ݹK�Z[I`v Z}_o>�cXF�0["���@��
1oO�3#*���Z�$<Lٹ	$�V����m��}*��.9J�85 4|O��d���	�(c�|m<�uj���Q�r	]1���!�D��4�P�&�Bjv�k<�a���/��1W�|KcV���@�����(p�By+:��W5ݷ���vF���/�G���`��3�]�-����L���OG�zd{�J��!]����W?KfS\q�|]֕��G�Q�=Y;�Q���nE��v;v(2��[_����ih,#]�5`p.3�,c�tjm9�u�m]�!f3$��֝L �c�2���k�@/��:�"~�8�*Dy�嗐��W=�y{G���.�4���I��Gn\�|�z@u��*��5kB8,������F$��Wo_�O�W�O���dK.��t��?��يwq,��^�p<&��5�E���%J�nRd�s�0Z7��f6&��Ƭ ����Aj�7�8I���g�@nm����ܿ4�_XۗY�f�5'��ЬPH8� +n�|5C���Ͼ�}��Ƌ�}g�Ե�I��\��|�+b���o�#z���'�������ӊS3%�!`A��7_`�� L��i�!y�Y��ZQ�~�#x7���d�5��!�������޾���ɘ�H4�����~Uy�����TҴ��㯭�}�c�NWk�=����n4�e���xQ�7�4p�W:���E'������:��z�%���k%�:�	�7;�RB'}"�'�ʨA?%c�ucm�<:�;���R���fu�`4��" 9;D�|b\�ؑ��?ʅ���_	!#� כ��Ih�>�D�Kq�e*�?�-�Y�y�HRD�����4����~�����3��5u�!W���u� O�o�]j�#�� F��Y��!h��<X����b�;���.�N������DS��_��凗�Ck�Bad*�.�5+���f��n�Ltʫ�4�Y	�h�f�:�C^*�h��xr�F�i��:�t�>��-ʬ��~YX�6З�m�̕7
a�i
�?��_���4%t��)��@3��/LO��	j9���4��G��p#�"!�=����r��Ԡ/q��+p���]V\�(N�}0<lc 쎔s�*,yܖ�Юu�w��}C�t^y��3t>�~�5'd���6����}�%�<��<��'fe>�a��w�)$.����n�Y���L5&��>�dA��Ѹ�'@�G������T�P�/��A�O���2UUJ�Q��N+�5�#��:��v@"�I�I��S �~������H� �O�2��JgR��`&5��Wb��E�E�o��"ZĶ�(�此A���i��T1�I�g����\�d��d�My�y���۰�&V�}l.O���~:Y��ǋ���@*Q.��"���z#�Z ��a#�T&ڹ����^/�l��fe�:��uۑ�
!?�X'j��N�!�FPt����n��.�� 	�z��X�9�����7�R���$��i_�4�v��:Y����@y<��mRm:RǠ��P�H>���ڬ����O��jX�:w�k�$j���Vٻ�L���U�I�OI��:h��K�c�R��	��Mpbfo%cch��$46Hg�3y�b��k�K{�ܣx��;�ہipuG�25,ǋkO�p�r�c�Zw�\V�C��=N�|9:�*�"t�|�>�����(�c XI������j���kl���q��GfY���qUAzi]к�Ӿ�@���X>"���sy�]�=�#4ۜ#��,���6�,�o2U6};����*X�Mw+!��#	�o�&c_��P@̈́�Wc�w��Q�B�7��"s�a�u�����_�u�0��H�~�ե8m,Gb���y��$o�+�%?	b6��l֜e���i膙9��x�<�?)u�u�T���= �-�XFb�VϷ�&��jS64\�J🻥�c<A�U��(L0�a�~��'`9ր��r�E#�ˆ0��Q�`3���fC�gCJW4���ӕd���t
�&r���'lѤ��� (Z��K���e�1)���T���>��4x�<�����s^�
 ���E��Bd��.��g��FLg�w�� 7���z�dY*9�dX��A�@F
�k��*��`�����F~��Rs(%�[7�	�2V<q��j��O�p�&�8��`=c���hŮ^\�ʜH���}����ܓ.fT�~�)/�����>3�-V�{@n� _,H��X!�S���K��/'n�O-L}I���[%���4>-k�oh�̵nn�Њ-��!��bHq��+��Ov��ȠX��v�w��;^��' g�_�ީ�IfiˉGܭ�-����M.p������JsYy��z���`J֙o����/ΊG&�܍���Ż��{Ȓ�%���ݩ�F���~���h��a�!�D��-{7d>�H�`nބ?-6�܃�.*"*��H4��->F������M�A3I�T&�K�9P�� E�?-7Avo��j�Ps�õhc��*�fY��W��b��nn��h���X(��	@͒�C>b�sN]ի;\�E��N�+�(#.`9�S���
���n�vL��#+���?=L/�F1�?�5	�h9��.�*�e�8����u��R n���[̲�P��bz#Y'�Y�+���uZU��{���-���n�k�,��c�M����ւ��m~촃��hx���NLU����z��#�1��EUUģ@NZ�jY~3����}���:���#���)��Q���$1�����@�A�L���o^IP ����s��Z�4�b ��vb"�y>Bo�(.+㪎�G��+�B����'��x�\��#���b�*@���*E��T��Ik\G���d�����nZ5Zo�i��'��9=��n��9��P�b@G�rl�������,7Q�R���.}��H~0S�o��c����m,�C��!�H�`�bڿ�S���_qxd6�j�X}]�l����T�`���S��C_�;5�a������s�ns �F�Jt�U����w<�Y��o��u��^���}̘�b��Y�z����2����s��#>�'y"(|k��������M/��x1Mύ���Gy�������Ur�Ųe���{���qw�k��$1�`r�xÕ������}��8��w~�A�2���T�N�~?$�
]���8Ҕ��B�i5Ց�����9�md`���04�pB �fG��Ǧ�H�؁��}�:���s�y�x
2<����� ��T�n����Z��?`B^|յ��1o�*�zd"�{T6�F\�{)X�[�!j������[�p(,>ힶP� ����(��"xF�Hj.���"L�	o�=FZ�=:���خ[~�L��6�!���CwY�����7:b�;z&��E�{�	&�R�wlhrQ]��,t��[���z���=��k�TW<��H�-����t��������	u���J�]��d@�D�^�ϰ�eU����,N�+?Œl�.�Ը�3Յ�7��(_�lw=31?�MB��
`~,���8��9(��)E���؁���\EC*|��0�*� ��p�YGdn�U/$a��l�3���.|;�����4`D~ݷ2A΃gE���^�pP���2:|Vpj�
�Z�=�Z,e���=^����+;C�h��6�[�h���(��g]gּ�C��hEw�%hƸ t�>�w��x[/��r��~%�m�I�fv�H�q�"�p�8}˾95ؘe�k�jJ�b�>4*�j 6-Zk�����g�L�`��/�ZN��ʼ'ՙ;��Vy{���X�Mϭc܅���Y��zHP9ݑ
�,A��l��XE����Sޭ]��=�/wR�E�[Gr?h�B5��2ߙ!-�#�k��Oy&��"0���e�݁w�O���5�Ϝ���m�� ����Ij�o�u�:)�I_���P�v�ZCg]Y�ʕ1�9rD�E��g���|������%�73G��ſ����������j�oO[�R��j��7�i^|�Y�c���6�
kt��2�e��g�.ZO���*׵D!��J)�Ȭ	���������,y���ᮍH�h.��=D�T�	NAs�'.�f���[�(e��KQI�ں[끈����N����,<�T͡�f<�ѥ�����ԫ�E.��v�5|��TU��̔K���� �e�|��jh����Lk��N�P߁k%���#.����#��φ�1%�
�4�;h���4��}�Ht4Fn�Hx�n$�����1���/�Ԃ/�7zU����������H����x�A���������CM��ڸ� E�3�~]y5��vZ-��#�Hq�L�_jgU��ϫ����&���2U܂'�Ql������LYB�w�r�����*RJ�;Â9|y���\��>Θr3(��(^ ��!T�l��z���U�tO�v���x7Fi�!��U�I����"ş�5<i_ٻ�:5��X�����k"W/EԮ���m��U����=�t��%hs~���@�R��uĬ���#�<�W�M��@���)������5=D	!d��q	�FE���+�"�}�u�Qu�6�(b�����W����{�<&@�����T�7{����M&��oX���\��
�������ψ�;T��ӈ�A;�L�cH"�&�/�J���7}�2��Žڡ����j倜�4�;�����cj�d��K3����Wk"ϧ�=��f2��3ۣ��E(��H����ŋ74����.�N>��z�5F�@�ж^�>2`kBPB����w��Wy�Ͷ)6:�1�-�`��[p�(���qJ�,M�oT�Z@n�PS:%/�o��n�o�$�_i���}\�Ҫ~!=�*��K��Ϩgk��3�����H)O��zhĝg���R1��[6\�c�ƷJ�6lr"�7�2K��HM�3�m� ��(���I8
j���N�����T4�It�Ŗm�����!�\�˺�@�{UUK�D�gC�8D+Y=U��������D����v"��
H�+��8(AH�5��>�3s��v��o��}(^��4l�T2��	���1�3��u> �C��R�;Qdv�Y=��.4}U�ٮ��Y]�п�4��Zg%n\>��p;�b�v�	�H���c\���\m,ە+_%t��q�� ���`�=}!Th���7��F�-KR��Y���N� ���ht��߿�vR�J���i���S��S>�T�[�ZV��M���0��2��b��I����உ���ѯx�+kuӕD�k479�7�
;�>Ǒ��E:�~����Z��6ِ��q�(�BѸ�cW�����AEplBR縅f�UL�~���)��S��f�qo^d�������M2B�q�?��6.'�%� ��,���n;����~�t��=�v�"����]rdp�c��U7�h�H�� �o����FOP�hXE]E?Ӟ] �Y���9T4�e�B���q�[��\�,̒`�;��SI����X��X;���.�19J6=� �̶E78�yB��YZ��>=�ҙW�Y�j�,��=1��ʠhNȯ�[.��#�|¹g�	�Km)���6�b��3�x�@���sy�&�����Cs2��E�m��r�جp����8��<`���I$T`�욠25&�Qj��$�L������T��D0F��/��r��D�_��o�@���c��������e�zFN1ւB�����w�eprƊ��uK iIw[τ�B�u���AE������P��;�,ܦԙ��/bj���R��0��n�򥽖_�Jq��S0-ލ����3�H$͒	`�t���7zq�Fv�$9`�J��"!��k��ho|���.V_�l���moV'R��g~_?A�Ij���Qn�6�Q�`#�(|�R��Z�z*3�����Ќ�W&����S��kv���傐��A�N置������!z��ЩJ��������6��?���ϕ&缚��w~y�d�i}b����j8ɶ��zx��3t4�fa�e��򼋝���.L�/�o��K�!���kE�(��6oڬ?�Y0^w�h�f�`�&�l�q���}�X�\Uf3Q5�̕������Om�`�8m��6<��Uh�����(\4�LG��)fyڕ���-�?$�,s��P�Ǝ{/
W��(��A_3"��t2���^�uI�-�dDi�*jR!��+a��?Ke����̘�3�Ab>d�Q��`ҥG��@��1�����\�(<�̣�����
&�w0��\{
0����)D_�
�t�5�'��#�Vx�)��(O\lSOl~S�����gg�%jo��V��Q��/�xBϕF�Vb]�����-��Fx�y(�"�E��Z���ȿ.����!e�\t����Xu�EK�;�-zȡW�9S@o��g|���p2��+yZ�pQ�"��#���CښV��X���k-����Ԁd�[0��!�ʀ %��*j�y{|��D��k�m��Rq���S����?��s�8G��Щ���S�Z�=���f�^�S�K�!���*�=�N�QL�y��@@N�d�a3�K{s�>9��]�8몘6;�>�yMr�{���K���U*�y��]癴�mȱl��()��}<�0gz�l�K^Ȥ3c}�rGy:nSޚ��c���MO�Fs�\�h,���D�ŭ�;�'\���\`�Z�u߶)�����X�N�)�K�JL�yx��Z	դ]����J9����䵋�fZ4�k$�I�/��ʵ)��pNGA����AJ�z�q:P��%:0�п��8�n!�|v��p����.�r��r�QH�z潻�tk�d�g�M>��Wʴ\ȾNc�|`���뙇�z�+@��EkhV���=���1��N�BŞ�8o�'�NJ����Ww6�yř#Uy��;��@���In���ЭR�*�q�=�(
�hX�>��&3P`*nW2!OiNH��e�;��7�@ 6����A@[C����-K��4+~�TVz�{(��@�n�f>���I�kx��/�&j1�ix�A�Ilm�Q��qڳ�ڋn�ڏ�����u-�j���L	v���u�=	��T�6�S�0?���l�u�%�4ե)��[>(��Q�]a�ߧ��oEuPD�
X��)TV�� �)��r3�Y����`�*=Y��,�'����0"�,�0�Xc)Y���﨎F7vbr��p )_f�w	����E�y�K�G]�H��- ��FL�����ͼ�^*�:�K<�g1�)'d��(J���K\v7<c�兊7[z�>O�b�'�����{��W�Χ��C3�XP�,fu�51����Ns�}�w��2�M��lH�ӓ��� !n���3�lR{q�C����bM�?���Z����F�b���SPN��5Px�k�����Qg�x�ܞIh�ļ5keGP��N��Ƕ.�u�š@�l��bd�dLA�.�R��h�eaWqKІ|��F-n�ﺴ�A%%�`�8����j�R�r�ǋ����QI�M4+?���f�:�_�����'lD}�&pѭ�7��aD���gg	.����1d��c�����5�l F N�Ay�zU량֔g?�[=��}��K.ϫfց�b̯��ޞuݘV!B7H_[���5�y���"u���x�ڏ ITH�O5���~���Q�*����C�#\�1�	Z���(�:r�p9\�LuP�jN?�ލ�Bj��9�|X{�a��5p��J�=�܏z���DP�$�����b0[�aS�|����>D�M��|���A�Z�ˤ �k�e��F��ucP�~�>L3M�@E�4����Cg��;����/�T7QR��-�;y	^�
���5oB��JCI(e}���G75�v�=/7M��=7��w����C&QP�iJNǆ���K, Mߍ���li��y%*�GS�C�#F-o�8d��$/�mu�)A��iV40�L:���8�r���-�l�Kb,��Lɘ�BN�>)��Jώ;���Z�
�Ih��ƋO��}�:��o�@rK�+"�>k'��r��̗�	�����Q���v{ǩ�{i(Qĥ��*�b�{���Po5��p�f�h�ц�e�}�;ز:�`	�����uJ3��ٱZ�伾�&���YԢυ	���Ȕ��E�����l�O~h�
��Iq>۸y�1/-k�Ӗ2
K����=�ð�[��- �Wd�bC\T_z���,�a}߶��߲%�cK>�	��B'i�dA���y +�������T61I�A\�$9�/^�5���W;����8*�N�2���dQ%�kG����0�5�p(��">��j#�k���� 
ak1��xy��b���і̥TL��P�k���IaG� ���d
X���[������ ���S�Co����Y�lP�?D�V0J�lxֱ�D�boE��=�,���F�%�߱��6�])�I��ʅ���dЖN�.��'G�p<2H�B_X8Mi��l?�ŞPс����M�;��?-H�&^���6!K�������X�O�Jg�߸�	~��z�/���9t������R���ЄW��'��LD	̳�/t�%���bZ�oѡEF����#(��	9�an�Z���׹�O���|R��͡	M*oj�����j%��7�@�:�後|�ǟ���$�>��f��L)R��,d�mU͍T�k�X��jJ�� V(�
#k:|/�s��W�5@��9�S�Ub�x�T���1m�P���pի�T�:D��ẆY�t��Y?l�m=SJ���/���_��d��4�v��ݳ��	�����H���0�����{tK�S���M9��kD~Ѳ�3msɪ㭠J�k�D��s</,�EcI6��kͨ�㒺|E���%����g:���/����әS�nޑ�x��}����2P�.��^���$-��ѵڝcm:T#H����;�ڦ��:��(j�E�ˣ��h�CU	T�IKA
�K~���t�� �
�,%�2���|G�������Ի�["�c����*Fe�>�@���5��Z?�NKܤ�Sv|f���p^l$K��Rߥ���(�,ͭ& �q&	��a����3���x/�ru�1�ʔ�m2P����T�R��F~*!��24Z<����}�83�eݲ�L��n�iV���X6^��G����DT��q�yX��ie�D�6v$�
�0��ۃ7c�ȍ�\�ik���u�+,��'�y�4��洈L�xE������.I�=,�O�q�Q{�g{20I�5X{��㲍��@���z)�wu0��3�Hn�m� h�^:1�Q}�1�x@?5�ćQ�{�*ovI\�1�t�(4�Y'�hA��}�1f���D�^Gwh���ߢ1�Q�y1޻��ژ�;�MT�/�-�>lRŰB���j�-���h���/|η���0�s��o�RmsT+�g�Co�Zl�0Z�{��Ӌ�CDO,ur��s׉=U<�f��\�]<˘[�����8�ga�
՘���	?��i]��J��6u�"��=�O7�5p�xA;҂74�o��PcE�N��	J��k��)��k�y��$g�G�eF��8B�sn��2��/?8��'Cjg��U>������Y9�؂G�%$��)?�.�S9&��J����=�S#��\#����T�}�ǘ6T�w�&7���_+���-��[)C��Z�3Y���^OJ\��ȵ�0�����e%���;)	R�ܞ��_&������CPaz�k�����p��h��Ψ��֚+��.$���@��R��1�ڴ	b��u�tu@"�˂�����i��1�l|��BX=^�H�TFqF�o�\����i>�HM������^�5q�SAi�x�7zӈ&?3�����Lxһ��Q~��8�r3���^5 �9��y.}�l���i�(�̲e��T��jZCN@�%ے��%ǯ�1�I0C����� DzK�;�J�Y��34r��<5�G�����w��m/;��3�E  [k:7�U���^R�������^�;.��ƕ�xU�Q��!Կ�"�&/�L�o�^��Wj#5x��O5
u�|����A8vpW�hU���8���)����|�N�Ŝ��;���o[��CNq8N�h�F���������r/6暑{I�$��ժG�����U���N��^�q�(=;6-AX��R�����N0qW4��ٙ��3UѪ&�FM3�yƹV�3��K�N�G�\y`(宫��Rp��\�MM��=�i��⷗���y@!,��#�ߍ8�4܅�72h^��%-�^����}�f��e�mej'n�>�Ao��m� 06Ĳ�l_���X�L��xe�t����5�ړmX��NYS䦀�"|�6_�y���^����8S����!ы]Q��'��`@Z�3���n!�?��������Lo2\^��BY}:�����oO�%%������_��J{��2��г� 4�\�/a'���Z��E�hD2ND%���T���V@Z[?�Kj��}�;e5�<J |�Lvf�̘GB8��:$����k��*�t�����M���Ӈ	�D�l��:�wd{y�jF��P��������FI���m�چ���n�Jrڛ3R_X-|j�� 8S�J՟���:��Ykd���	�6�ͷeMVFf�S/W9���i�6�h
�"K��QHe�7�b:�5i�q{c�փ	+^�̞3L.�k�!�#A�cb�Ռ�̦�x����ʺh��΢����x�t;M2�(��#jb���5��)�Ht��j��)��H�.�緄gA�~�Oߏ��f#E��P�+2�2��l�Ǜ��w����W#�O.��@�osE��r��	`{�f�o��?P�Lzo��`��s-8$Ҧ[+4�d�I�U��Y<��u-�{X���o�?lNv�O!��uj��K��g�h,�&L��D�BN�u�X���U�:V�}~PW�m2[|$h����|�=D]uPu�178�$�5 U�Z�m��U�5�.U@��<�ij���QF��}�`��"�2�Ӹ*�@{�+]0R<ZH�{U��0I�G��*�9߇��o`������](�@�E�{
�"Dt�c:d����A�q�J�m(d	��_\|�qT)�U�H�T��HW��{���>un����Ak1]���ڝؖ�t�|OK�����Ժ���6�	�;pХ�V��Rs?l��#��|��w��r����4��S Dn����Ar��i��m�oGت���&���;C`rg����z�D󇶧��C�����A�S���3Jo�Զ��1����r%�&����g�~kD��A��Ps�
��}2���E5|o9?
)�n��J�+���&@GJ�8����K��� !�f�U�'�G��*����;�!�y��å�LC�[-u��-�?������Z�;�R~PLz��aZ�~�1�@�u��=&�P�*�=��<�,N���G>�>s���,��x��z!Xvb����*����q�
��^����U�=���rE�_<d��n>+�^�w�r2�&�-_OjB0��rlףG<IE�qqNjp�����-Iٗ.��Ҭ�U�%~X��ꛊ���o|�����N�����y6w�(�������i������p�2v�wv&��lj�~s3�����ƅ�ZqHIq��xL�x���ރX�&YG������&��x|��颋/W
T�L��[��jHJ��2�4��p���I��h�*�H���>�C�J=tgQ{c7���2} j�'��X5wWv7v�����@�ߍ���f�r���L�.���)dPO�mǂ��*Ԯ���`?M�x��iH�t�V�m��t�:,�#c��� ���N{���m]�\�����d mʟw\�ˏ���=<����*�����gb�nc(Z�Gr�X"��ډ�"g�9����T�9�!o1��}��Tre�D3�P*��G�㻀�Ei�{�7К���|$����A�:�����Ѝ�`A�Q{D��qm.Uİ\@x:	2q�wf{PR���������ԼV՟��/L���E6�a3�O4)���9u��}7�u��г�,,|z<�%��``콎/���[���1W��F���x�|�IR7y�狚J N{��N�(x��gu�f^�z�ׄ`}4��P�49�����8$���4 ����E�,u��e�LM'����B��΍h(�Ř��%a{�E��s���8�/�T�-��4�u�5mw[I�S�CKhm�w��p�0�4łLvv���S5�|�(���J
fV��.�4�|�D��e��>̘��e��愼ߟ��L���8� F�۴+=�6�΅�@R��lr%�4��g��f�{ș<��D���_��W}/��~�L�xj�_�(ڶ�DU��띏nvȤF"k���5�m�kc��7�r�/�W��iJ;����������4��4"Ԉ�a�^��t����t}�Z���nUW��*�m�Q�(�)ԗ�J	����l��v#l-�M�|X�� ��ck ؈Q�(��A5`r _PI�L�/��T�d�Q"٧"��I�{ʣ�fF&ZK8�åQ�1�$�|h�϶�ܚʷ��.�~��WkX~�m���v�xғ������Q��/t���Vp����w*`�~�y��i��0eN?����̲Uo-H�Nޥ���&>���ptR��,�2�`�t�}����<0�`�D|�pV�i�J�_��!����g9~hq2�cNT{Mk7&4)�l�����U�\A���<�i��w�̑.'��x��w���S��#_�u Ws>�_�g&Yx6,	�K��9��*1���ކ���=����gq5����G���`�1&큼 �I�o�j���d�Sy�B�76Qg<uU0ܼo 3-P`ރ_R~��}V�s�L?�ғ��̧�P់!<���s5���7��
�5:�;�L�yc!�9̈́+�eA}p[�Q�-�b�v@��F���o�C�����L�-.ו��'�u�=����{4J��������vڢ�9��+t-˦ԏ�f�zN߹�tQ[!� ]ͯ/��S=��x���q$']��9�U�q�쇡t�)`2�r$�Yl6�=M�\���Y�KV#A�O@R���mϓ��]`���q��j���Y)pᆠ3)Y�$�P�2t��=�Q垱�����<��p9:��)���M���f��hC�vCm=�T���+��yN��������u\V%��� ��LԚ���+�f��?�!?�9��
o��EK��=O���@�o���ᗐ;�&>�&{�F�Ŵ�@��b�(�>�&����$E��˰9d�̛=op���F��IL;�d���Y˟���A���M����a����<�����뻆��o}(o2N���E�fCb���jN��q}�S�uhcXQ�M$�aP��8����?�֥;PD��z\&(�6v/h���f��+£넃�v�O9"��}����x�*ܜ3��G�-�m�1��TY<��.�<��sQh���L�
nW)M�� z�UvM�=ʺ�"�� �i# IX�xL�q"�wN��� �j-��!��GhM��U��6�ꁟ��lI8�������1">��\
�A�h�]�kv��˩��Y��([r�x�)��ﳷ);9�b���W����Us���bʔNT4ç��
�]����"q�Oۮ^Ո�O�j)Ҙu��D��� ��$������J^�I�=���`�sQ�����A2�o���"�������3ok5nͨ���T�	+�������k��@�6���<��?�͎��G�>%�z):�7�?c�36�9J��xP�
���\V���@���_��p{��2/����٤�I%�zmn+��sc�/[K�����(g� �?�W�!=!9�I����w�ˤ�B8�w2��f�y`V"�:�M��/�&zP*��E�]%Y[�*�nQ��Dڹ܄ܦ��ڕ�^au�]o\
�Աr?��e��*Maq^v&Q�,����a��@_~�U�ǽs"�w�4O���=���!*
!�t.x%}`�.V��`A�
�h!jb,7Ԛ�(��;�A�:��ap:�:r�T��ZK��j����h�X��̪���< ���xi��r�B����W�P��"���4��(�m� � �)�GK�n�^�P_qL#�S=���oL0C��>�'�c��)�96p$����S��r<�K^�>�Pc���Z���p�G3tl�4���s����P{5up�1�e�T�S���t͊�c��
2K	w:�U2�"��0�ժ��6���{�V6S7��F�7�lr#OG,�Zq#�/'�S��"
�y�Lk���q�28���џ����h�c��װv!�eK[3��Ty���L�� ����%�Q��+r��1#�B߉y��U�n��8����|��\P���V��y�����SXIצbȚw�:���L�I3�}@�㥱m՚9�["�A�RS����SGU�MP��'���
J_�+��b�+F���<^Z���pS��D���+K�����F��e.3���z��\sPJu��7�C�Y�2X�1�X�SJ��+٭&4`^J����o��<�[Jv����P"֛�'i�>,eXE-�~�Ç&�į���E�-��N)@��s��(_+��S�7)-G�QŌv!�"Gr"s�)����� g_���T�^]ZH�����Ŋ ���<+�~���3ѯ���o��,�{��D|�@��J�����W~��xN%��**����^���\6�&3�=GF%�tz&HE�����{_aJ�D�r)�����X5���`��
�.�LgG�����~��),m��'��G��J��^�~ڈTL/WKб�
9"�������dx��N�Bn2���i��+N���e�;��D%#k� �3,������d��-hf��E��o�C���-kV#v�������ń�v��_�g$��	�,߫8r1�/]'T��!z�d��7�!���3��[9�l&���I� �.T���Tԥ��ڂ|����6N�]t�������s��ȷ�C47�A����~oH;��A���-%�Lj��`^9b��.3��R�2�	����hZ3���H��2yR8ԡ~��R�\��
=����]J����3}�c�6�a6.�SG_)�$��1}$���5��8hV�[���cܞT�_l0�2d�f
D%�
�������	^lZ��^\�I�I���yq��P��x�4e�ލ]r���X�j�,���.��yN��i��B �HF3X�����X�����B�0�)��x7{�1k),`�1��@�uv��D`�-ླྀ�>&`���1UѦ`���K:	�o�tj��)cС�JB�;O����O1�y@�D$�A��t��_�Cݒk���9�:�QS|&�|�� �>Sl�K�w~�&pn��-E �0<�
)���{|Ǉ���_��K�wf�UZ�eg��%�]G��
v�����x�q0ЩaG~=S��T-C�S�M����+�<L�׍L��VI���5#���)5&~��ʚ,[��D�t�DL��0O�����GC�a�����'�
�N4���t�jN\��v��j	�����M���(�[�Ǖ��������{��e*投#up︆ZXI��[�Z�ؓ=W�q�-��"��n.�Ks8�}[��]��k�7�R��?Z!�ȭ�
�n�#b���J�?<���M̗����nt�O�2�@V$�7a�~t�1͌�1g����C���:�@��� [d���%���K�J�(xk~~�Ʃ]G�y�(R~A�c�� 8r@%�5�»\���S�Wq>-��NB��CH����?�`g�*���Y���EKrΓTS�A�krn�w�P�9^�Lv~!3��3YP��ɺ�a�~����J�D���<�J�}w9��{%,��>(MH�
�ś�:���������4k�Π��Hn��I���]� ��<t]M���۾jN���*������͊����&��2(k7l>��^Po���a����Y��΀��c�- ��o8X�g�Z̖Q��GuOޥ�d ��p�9^��׃F�����,�A'�e�)��Bi��ݍ�I�*�.4D���p�\�H���h`��=��,2��F��8�_ڀ_����8�v�C���ܔe���7w6;��X�[xʛB>f��$��dx����&Q��u91܁�s#�s�6Tor����+2Ǧ�8.� �=?��N6�K���89���_e8"M0C�Gq�ڪtxN(��ش���kɗ����9�-0����#���<CR�L8�ՙI�>0I�K䬓�I�[��5��� ��O�6����
��҈|5B�
�b~;+�c�3G��vE]��"�7�g��莬T�jL���!,��i2�Ew�&�T�c��U��`�/�w�t�rb^�L|�׊��m���2χ>�,s.���<3V��Z���l�m�1��(tu�8jd%��Q��I��鸑>ǉл8����Vm�5�t I��N��+�P6����&��*�x��sr����{��}�i�eO}��ui1��
��ǂ�K7� �����ٛQt����{����������J�}r��k����_����UyJ~F���0�~'����ԁ+,�ᔼ���n�x�ݜ��A)��;驷����f�=� L�A�Fec|6���1=����԰X}]��W.��0K�����Q�U�;�/��I�}�ل#a��+]� �����L���L�x:�q���t�n���:p��Z���*T�P/��7+%�ǡ�{������i�h��V�6/�X[	��E<�`͝�H�OK�ӛb���x��ڈ]8�iL�G�����!2����҈JNA4x6�ƪ�Z��񧍙��l�LE?��CQoO�n`�Sr��p	D����=����{j������rW�I���V��-$l�i�P�Cl
���~�o*iW�L�d�`���(:����D�4;�vyY�,=}n�k�w�������`K���Ԃ?{������c�V�8;�Nhz�{P�"��Ŋ� �wm>�-�*�=I��Y#u6��T���K�+���r�\�r|vަ����ױ�C���v����e8��C�h���sV轫�}`օ�h"�:��G\��5Z�և�&��]G��1�p�J�|	z6������Ч<ހlhbؔS��߸�d`71��Z��=r4���_ڧ�3戜��H�K��U��/��]�LL�㋜���}H�j+aϹ����>T"�����)�*Cq���#�ኌh�	9³����Ћ�n*��nVG��,��IX?�\�|�KE�B�EYQdf'3`�3��G�"��7������#��o���$w*��"��dg�����#r�A$/뀪�R�]��7�o�+�c�:S�T��<��v�7C��F�X֮�7J�`�x����4�����sI-_�ăRDb��\���d�a�,�j�˥X]�IJ�6c}�}�Ee�嚙#	B�P�pR~\�z��cE��ri� ���3��$�˙raԴv1��rd<V���%a-]&�r2�,IQB���� ]��%��G	UCcM��ͩ�i����p���N�ۃ������j�"�k��
���������T�i�y��u^�Ύ,�Ӆ'�:^�$�b���E�|0�'yiL���<�m��Ǉ%�MSA�'Ʃ��I�
&j��T
<�>�w�Q	�}C���yΫ������R���2�CS�y���<A��(n����y3�̦+@�_���(6`��L���ȩ��A(.���w$1�$k���r�����
}Ɯ������R���)_+5��!Y����@Q��0�d�4��H�ڸ�v-:�utwj�h��:��79����f��LZ�$ђ��W[3�Bv#���X��
�{��>��G^k)
��Pm�n��:cY��Ze�$WҺ�����kձ�x�f[�a���Ѐ��n}g�MA�ؑ���q��[�84�`�x�Q�(�I��ה�g��q�9���[��|�Щ��Ðx:4;i.�й9m&��Đg���;��/�E���H絜�u5�a��[���j�Ed���6#�XZ�#j�+����-m�����tV�^B�T��W��-E�$�U�>M	c����X��T�zя<�)ʷ��h��"�``{B�렢 ��@Uw�t�B�����e��:h �������W$4���݁��U��r �6��X��R�e�'���)]��ٔ%�g��K�)..���E݇�{�f���$r	9�w#6����×�kh�Ձ'���G�=�oj��xH�t�[��������)��Ŝ�Z�{���M4�ؖw�l@w�#���c�qqQ��y�6����93�������r�>1DN3]��4��N}��g������X�X����������*�ޗ����� q3�T��(<��{���=����sn���z���^�L��A���4쫄���t�|B�Ki�i��N|���ё�RC�%�g�e�#Ixn��iW�Nb4Se�<��d��-%�1,�߳j�Q���a�/�'F�a������w:xKB���D��C��k��d恬�@����d;�oU
�'��!3^_l�52mN2o�`�L�qQC� �4�C<=���k�2��(w3��A��Q���D�J��H�23jػ��$��[�;��*S�^��N1�V���U����lz�r��p?P��Z�����>�x�𴠯��P91=.S؎J\��f��dK��-e�lfD}@�B9j���)ZN�����o�4�W#o�:�����~���bօ�dW+��䗃m��*��J�+�gb��79D�ma�Ne��b���;L*��)�-\���I��߳�X��^#Q��$�dO�խ��	���es!>����A�j����� ��{Q���'��20"�|��5 ��eG9.���	�O
;U�@��Lzi��?��:�*s���Z����_ⰴ��L�����ͯ���g�/�+����u�����������}���'"A�
�z6��Vk/lC�Zѻ*�Vu�4(%~]�f�.l��K�) ���75�V7\��^��s�;�B�/۲�#9�C�E���	n.��o����@��G��
Z��j�Q�"�G��;C=��. �勐���L& �2�kmw�N�!���3��Σ�E"��VLW�`\��ėUX�<�CN�%Z<��r�@��|��k&�nǢZm�n*pK��ڽ���>��Mս��j��&p��3'fCs��*�߭�a�y$�����/��|�=xCw��CD�qn@�F�G��x_�A�r/��9�eY"�����PA
vY��߿Q�I'Q��`�O�2�U��[���?��ϸ�/ ���k�fwqf�)3:c�q��9���v�	��� �p�W]�b�X�\��<.O_,p�z���TiqC����Ԑ˩wї����Ӆ��ͅ�K�T|*OC��0Zֵyy<����������M�xޘ+r3t��AW@�-?���Dג�
PaOh��\��5Z�E�#��ߢ�!�����i�ne��x �Ҷp�2��z��}jc�Z��Q�-�r���W#�y  7�L~��c�l���'^(�޸	\3�[���M��y�ܥ~�}&�����B�t�o�-29 �r�4A�*��6�f�%h�/='�oI���8J�Y��:JC��b�����4�L�c�C�ܜT:�p7P 2?������z:���-{����vD2Ja�F��ҍI*���D��n���V(����pu�U�ssk�"P�o�E���hI�.�p���^��Ht�?~B� oe ux���٠��qY��]��P�Y�zˊ�Nxr�
�⧝��X-��Ӥ6��K�ׅ��푆��f!�ɲ|?P���<��chԭ#��Ъ=,��
'N�]xhk����Ď�s�o�6�(a�ip��w������
�.[nI��%A}�����_xS�6o�D���0��tE�;ϡfU�3P�>�{e�-kj(~[l V�����jCN���э��huw)]�Ӕ���An�h�&�9W�n��=��v��]��(���)�=,�+�n]����423��(=:�R	���6��=%'�d4h����O�qd<����r�NU\j����fO"����"���O�A����`��Y.6�b ��7��d��􌴞�r+��J��7�[�������R�\���,ʨ[O��6!(�)_
2e�Zr5����c���TzL0���X��,F)�p�i����e��I���C=4�m�Z�$�GӒG�G#�@l3�m�)����V��n�3�P.��#��_���y��\k�#�WS�Μ���#�#�2蟧$��9���Hႚ��A��r�1�#�R���y�k"J�#&����3vg޳t��_tzݸ�ڃK���P��%!�q�~���j�g:��9!��P�Y���$�k�~���H�I�����^��.QJګ���Ma�B�e����Z6펇�@��%�8�i��T��X�d��ϩA��yb6����9���t�Opj~0e�f#�7�SN�y���I�Y;ǉ�Ze4�
����^����3g�c�p�}�c؊�va\��9Xi� R��qј�v��VJ7�l��'�Bd�!:-�c}��i�P3Y�	o.bn�д��ur���9�s�հ��`?�.k������yX���x�0uOSng�,�nf�q�Mr��?Ⱦ�#�.]��c�x�<Ed'uP��	t(���"p�;]R2��&Δ��bT����e�|�SD��;́�tL��Wdw�[��S+s����.������+�/3)�(�����E3m@��N
C!/�L�Jw
ɷ�[r`�G�:W�(� �������F�\ :�p)9S���3;��I�{ʒqgK��D������"����- $���+��+�M]��0��	�e��]�o#1�9����WSu@�n���Q^4�˹�=g�r�M`p�:j�b�JͿ̂�$�sю��OL�B�}���d_;��&��2(���n���V�Lں�C@'�}�1Ნ��Z;����p;ڥ%l�d4����	."�U�1��C�j�v�����h�9�
��z۱K�Aa���,���n�B�<��Z�V�#dh���V����L�+Ar�<��@�B�^�������-�B[�J�;w>�/�|�u7%(�
��O<���w�b�!�j���`b�a�!���ȅ�ȇ�T{bMY@ˣ�/�Wcl���[�^P�N?B�M[���7Vn�Q'��M��>j�o5F(���ȗ�ڹ��>Zn~q^����Nh��������Ѭa|�-q?M����>�K=�|���h�C�Zp.(v9���i�:`V9"��$N�C�&��Xm�ױ'�ìR�Rʊ�ޤ���44"�X����8)6[�YA��/�O�q�)�m�䳋�?��F�{����B�퍾�Rz�La�*Y�F���������/���7�(�U����\��L�YqW�ĹW�ϸO�)<(���0������`l=�H
���åb��tmc�k&���.(�<J2�����|��r��h9�&�lSt�b�SLw��cΓ0 *����8���Eu!��4��|��q��)|���v'i
W�2Q?�M'o��o�h\���<�l�[�` � ~)�^6��"�|�N�`(�8KO��$�՘�����$1f'Q��m�Ј5ĭJ$X2���}+���Y��+�Nqfj� 	���_v��dV��4�����a�.�涰^5��C���Lb�L��]�C�Zx�$�mŪ�:�H�g�+EI؁ć��J�P��#e��	R��
:���x��o����"�XU�Â]��̭�u��ZN�cX"�cv����]k�<wt_�2���=�7�D�:` �}�����R�OE@WA�`�`�'ԡqQT
���D�g��Oc{��CPvG-������ܩ���G�����^?X�;c���Ɵ$:�e�@PAh�܄��s��'��X0"�5 !���G�Zr'�A�Ɨ,a1�Lnӓr��2��"����=[� �W��^�H|+ �ˣ]�GV	,�FUJ��a<�ӣmA�_�3�5z[�M��So@[��`���s�%���mZ�����^�W����X5�T��6R�QH.����5];�h����,Y'�K�%�=�
�V�Y@��1x�}�f���c��b���aP�����oJ�:-�߸��eo��:!���g��ұ�WL%�<���U�312��i๮\A�c���\�� �D;Lf�WĤw�o���+}������.t���Y��O�#p���1���W���Fa���+�E��{�Q'�\�lN�����X�pYcc�hF�����⮿�UԲ; _h�,�A2)�E��{I����~Vv�N��x���d9��Y��r�4@��2']i�񲬥������1�F$	��������m�HK*����`�'�Q�:��ѳ��vZ�7���D�JN��=[�-�.l3�e�6rB�!圪a��i<�'R���b���]
�|�I��?��b�%����@T�3Yθ�$!���>��Z¿�ҡn�����-�jM���[a�:��n�<����e��30۳��נ��V�l_ӫw�<����5���L�g��E���a/s£�
JB�5���/�L�=G����	��]*�M}jy��Dڣ���N���gP�5Tq��hğ7�m�c�~�(te�a�l�]�*�(@�!8m�6���d;S����_��[�)l�����f��zN�c�,��������VQ��T�F��DPs����e���kypMl���S9#����KX~/�����f����6�ZW4����i��M�
�Õ)7����썤�%��tk�x�ۈ�ӯ�w�	l���O���8����ƀ��``��n�3`Fh���p;�����'�S3���/_ �����t���
�8�m�-ww-6;Ԩ��ތ������<	F�����t�X�? ����~�@�leyb��'Ԅ�1�h���w��7���a���aV�D�*�pT ���@/L�~��l2gEC6�r��Qe3��D��<n'�%5������4�[��$�R�使^�k�� �vDl���k�Js|��F��GW*�+�*ү�{cN��	j�4�?V�@��{雁����V�	ٵ��^��l&��pi�R�PI3n����ߵ�J�l5��3���Ơ<���sC)���ʖ�<�$�QסR����J������bɄ�j�)���'�7ч�1yO5������θ�bĤH)R�a&R��O9��M�x�hŃl�[�PU$��TA�����T�{]i&���1�J@�hV:��h0�y1�q��Ƣ*^C�(��c�N��U`.���pjwl�)X����x����g�*CH�X� �Vk��S���13�S�X�L�b�\����uk����p�1���ZJ?�_��A���v�K���R����{��$�+؝<�����1���w��j���Yf��"{l*:Ӝ&
%��@��
)9��j����fb�D��݉Vl��!�ۗ0�+C�6����U�"��S�kZ�A��U3�-��ޚ�H���8R�����mv��q��+����hH�(|�˗�l��?�U�j1b��>��p��\���aW�C)���� �?�]�=�����0��`���(X�|�w,eW�>m������\�Ot3G�t��)�ћÝV �S��p��	� L���q�Rev��������f����K�k\�~��A��{3�D������D����h,.z���1v��v���w�w7��'G��?�@(W��j�ͳE�CT���QƦ}�Q������
�j���)�ۦ^hh�`�W��%��,�y��ٚ��W�w,	#;���X�
���j��������d����,�=��e�Â��%�QsE�EN���AMJ�M:���/o�j�g�5q~�ńN^���.����d4�P�o�n4�Q	�q�v؝�o�N=�Z�z?N7�N�[���W�;+5�u�2g;c%�2�*@�����q���x2����Q��G�2~�)����<ͯ���I⣱����M��O����J$�$��D�z>���xP�q��6 �aՓX����x+ #ܸ3@P���e��p����8zZ*L�-�Z�&��S�^�$@V�������Ӿ�F��S��8_'=֑�P�	-��r� ��9�˗ѥw��g[&��?u�d���T����봁�����;7��B�-0	�>�Lxʢ�0���V��z�)-H��a�s��k����l�������v���D7>Ow�{Df���s�#�	�������nt��i���i��Qm����o�����Z����؞Z�]Z�A��C˷jJo�<V7�?x����'
2��B&z��a��Λ��	F����%JxQ�X�|�����3N�G�˅��=�����)>r����yl�F���BrP�.]���3��\5Bf��r|Z���=>�l�AUZh��O"-�ɪy�����4J�m4�#Kd�B	����k���'��󉂷<��	�z59���"X�I�S�j���nV��H/�)৊݇�OU>f�
1������T��s���3�Ktd�|����'wH4��E5i���уEE�$ִ�D��g�:���+�H�͔�X(�I���\q�)�_؅D,Y%r�y�5�<��[O�9p~B���V�1a��Tw�\*�~�񯥏���'�,O�v\��V�q��6�X��L���k��`[[)lj�As�y���X/��Q�*k�����zM���<��M�[��Wi���$�����~|3΄fC����6��-`�Ƀ��V�i��֢n�G࠘}�_I8�g�WFc3���+q�@#���F0���U^5Q�{�h!%=�I�i�����m�u|��/�kz� e�[���{����,����p�g$}�Se9�Pf!݁�!>��hX���?d���W=�j��ލ���	;C7�Hjg	GC�>>�POZv��ݭ�l�@~� ����R~|�WI�����0g�R3�����c������J���FkFۺ��"	��R����h���j�o;j�Em���Y����_��c.lƿ�XK<i(� �<�
�Ԏ���ҘE-Λ��V'gOy��S.�SP��5�sD`G p�{V�zhsùx��,;8M'�-G�OA��I�Ә+$'�s��$x7� 4δ�=R��~8[`o��:�*�{T��l�,*�����J(�� �ʞ�tE�Im���kwp!���R`�7��%|�	�-���Փ2;����laZ��|�o��q~e$Ge�Ϊ����k �Q\����((I�l̉:������6��.�P
���.m��M���c�ﯓ��� ����Z�`���B����b�Ŧ�������XI~!�Z�_"p���qq�e�#.or�|v�CەD�+j�y�[�i}^d�T_�J�+0 �{��O�t�-���?|IL���u{�+[E�Q]�m6AH����9�8���пk]n�<82� �ԣ�D4��?��WE)����Fnt&�ұ#n:�� º���W�L���)�8�Ru������p�B8��cF���7c0h�'��>�	x#<����g}Uع�v� �u9����HӀ��+���=�J�M6�ʯ�J��S����m*�v�����ޮ:sL������U�V@R�ڬ�����&��+����>��P-�H�ǋ~��_��>WKOڵ���(���?x���U4�W:������;/�>�����˵���o���F�}`��.�Wܘ|ᡟ����DX&�'�p�AX͐7�$��GU�W�&n�R�o�0��{oBÐ���;�^5�)��h^ý��G� ��0��{��$ѹ�?\|�ŋk�d�Bk^�!m��Mi�����j�B���R���YV��{�s@������V�^$W�1����h�8����qA��||n#DN �K�����5] L�����ҵЖ����d���IʮdQ���!Qiй�P���)_HH���s����HF�\eS���H��6c'ju�z6�o�<dH��6ae�OwM��8{�������8���
�ꘅ�byO|�[c��eE?*��N�,�	�K�W�j,��l��S�IR�ʶ�m�^n��e��5c��(�vO�J?�ֵ!�B�{R::�um!�C���ߓEr�����7[<N-h�ƝzR��������x�F
T��Q�Lb��鰮�G�F���0���5�RG�MwqE��sT#���]Ha������E���Y�� �����#�#䞒 ��&�Ճ~���@���V]�o̤р]�>�Plԇ�.�,��E�n% ��k�xC��Pgx�,�\� �7�@Ln�#Pfh�4ٓ�G����}	�*��w{v��g�ò���t����_��Ǜ�\X]c���b�׹F�^xlC:�'�yrc���� �F��X�6Ԁ�d#�4�#ሔ��±Sq�E���w���'�5O_����t�T�*v[��:�J���0ҹ�dT���l�%��D�:U�{kE�K� ,���Pq���?ݡͪ;!>�|k�:��Y�'i��Ul3��w{�4i��c��,��Η�-]���UnY���k����e�x㥝#��Ј)���.������%��g�~`��X�Ӥuh�9y��<+����怸�(�pnI��I�����@�OP�l�15��E���,��;J����*p{bJ@���:��\�}���m٬V�����N9�̢#?�~3�q��Ep�(��r����j��� �f����ݾ3���nl��+R-�x(���s�����ʹE�<�fo���or�)8z�6+;!�����$�0Eq�7�Q~�-�W z߭,���+����h����f�x�nv��V��6���֖�z�`���kv �\��1��`�r�,��X+NS7�S�a�,=��(���Z�Ɣ*�ע���(p����Vo�C9�Y3�J�|K�4u"
d�@��+�2�F�AwY'�rH��ي�z�G�&���`B0fca�)X� 6��iV��_8�`���!���z4�YN��|��ք0[N�'���4��X��1b%t�����*tn�����v9��H�bC�6N��� D�
�P鱉���z�ҿ$�!���#�CR��w�\p����Ȉi���X%l%�K���R�s7�c,a���r<IgBK�s��ԕC��ߞ�8��o��s����"?cƈׁ��7����|�yc���M�"^P��p�l��Aƅ�W��6���o�C!N�	��5m7g��om�d`�c���x�m�H�HW.�I���$��~�?�m���=Qw���<�1��*�T�	^����){
�y�T���7e\���'O���o��^C��8��е`7D8��[��B:i�C�@�����E�(��K=�m�'�����k�����x�*�e�ЧK��j�-Ʈ1�Qe"�f!0NB�r�t�^k.��FL�Z�x�v�^%�d�
�1�:!0Y�-^b#Hn䡼1PL���T��}�,d�k��nN�,�ׅ�)������,ûB	>�32�_�!��2j�6D����!f�K��0h���UŠ�hI���,�c��`����U[���AX���!�;��C����ܱ]c��7���Tv2�e-��+Y���8���RR��DA%mmz�6��g0MQ��������o��#��X����xς����|�:ѵR���j/��[O�A��������y���E�1���=eN�%�3FFq�l�2ձ�?�|E�:���D�G��P�
��O$/s,����oA1�hN�_�8w��E��E�<_#�����©��	`��l�J��_!EX�]�s�Y���������}�p�*�2*�Z,R�����Iٴ��bjm4�����O�f�8�Ԏ�+P�	�ɧ� ���&/��^R�M��O7$"�m/��̃_�A�Vp�yV�pK�9���qSNbCB�)̂�j�g����_�_}>.��43N��NK3%K���-�^���k6+viR$���<��]�����]ي�)��ݼ"�5�b=0�e&�r_ Kv��܇�IS��<j�4��8�R
<��%!r�Ď�H��k�1�y *��t\�	m���k4�_�����v�+��(ٳ��މ�Sn�	!w��}�����������4���/���g�i!aeԧ�UN����� ������ɹ��.�8M�/4{<�$�p�w�ύ�'m�͑P�Q�[I�K�Nz)�ͱ�����e�0P18J���8����c����ӄ���'�&HB������_#�ܚ=�8#�Y�М��3��������6�qfh�0���p"�����'�+B������r�ġ���nCrG����M�g��ɅH�C�yc�pܴ�h-�J
gV=&=pV͂�L��m����#L1 y���Uї|���l�zk��I�f���+��C�#�>����7��ű�P������ꢱ}�Y%* �c�2�~m�PL�؆��Pf[�>ɟ��&�OB�Ƙ�ݶ�Ҭ\3C�9@�h�ǒ��\��S�=5G��y�C*Q2���/,/�~�é~��D5Ud]��Bm�AD�j��օ�������x�<|��IPWpGec0�
?*$j�J�[∆.�Z?�8zu�!���I
^0�A�L�mu;[��+�T
�l��Ԛ�@ghJ@�L��z��@J.�Kط1�?���tѻM����	%��6�8h�ٶ�W�'�-�THP��ܺ�ˀa1bW9��E]x��z�X㐰������ƥ��[�m.����N�9�J햯CG�=��ͧYu�o�3�Lʫ*'�]�~��v��*�(���Nm�/�H�2�L�m,�:vy(`�.ۜ��iǓ�=��'h������pXh�ư�xﱤ�)���y����ے6V�4��َ)�1�G�[��J�M^u�6F��n�_g�"٭� ��rGh��"�Q`RJ��LvG(I�%�l~l߯J�6�J��{�w�05r�e"`�cWӆᇘ��r�'5h���>���hOc�Hi-�n ���bV�Taz��g��TX�J�M���h/K}�	�z���eD����l��d��B$*KY�ݫ����4�dD}ia�
��|&%��w�����k��g��3ӣ&$�nM#ґ6�8�X]�O��3��E���o������<��ɢ�h������)�P��*�(�`�"��&�Lia=«%��;��؂G����F�`���,l��*����ь}sH�Hm����,ߌ���g����' j�Jխ`N"�x�6����j�t(�'�����9L�"'��r���)�D��L�����aL&�����ٲ�3�̪æck´.���_B�}֞*8älV��֚��˅!r�%�θ�$Ī��xH1Jo³<�;Bj�.�>=N�յ��#��� ����GeA��qާˈ0�E�u�-����%�V�R�l�,�p�$�EM̏ς�}�!ꍗ�?[ָ�D5�(K�4����Ma���@��:D�O���t;:db7���_���Si��,CN�7B��?�0NQ�ת�mj����!n�-���Gwg|�����_����ݍ�ämT,unpr.w�=9�ɬ-�HuR�Mj�0���b_a��|�ׅo�N�?rTY���iLj>y�q�<B/�8���b��rL"Fy�no7�(C�w��9�a�C^q�c��@�%��)��1��K��A��e=%ToLb5�L���w.�.��!߸H�\����p���J\�V�T���7�(��폶ɿ3�!��/�n��a�q��=���NI�M�,v�$��Nie.cf����~�żq�q�YE[���m���`���Xk�#�t�x)�en�^�e�����*����q���xXk�����Ґ+<�v �$K(�����_'x�+��[t�	���|-���,��A����'��v0����}��Q��U)͘w���\�u�|��o�e;D��(��o6N��t�͝jb'/���g�Ezw�m8U�v^��u�a92]8T�H���R��7Gnz�j�M�m�� ���/Q���P3��� �Iq)(-�����{���)��UM����wM�bHaT�!��jCG�P���մ->�F-�Գ;W����Bl�ò���F���J��v���k��]����EL�a�+��\���s ����fzT�u9�v~�`9�[1��O��U7�&`q`�}lA
�w�u��q�p�j�`U���4��d�4���U���w��(k�8�����ֶ���a���T�2�++,P+��6�.�?��q��fTM�~?����5Z�Ma�F�����/@<E��챍LcfI����5��,7�hm��_���dxq�l�IkJ-~0d�_{�X��v���[w6��?��cu�(��$h��i�S֙�0��@5��'.�_�b	M"���y,�<5��u��y��J%�,���.��W���*u�@#r�Hw̢iJ��-�d�-��
���k����;�AVu��I�)b)�[�3���K1x}<�z�=��ʰ ����՝���D�@ѷ�t�K�T�����n�9�.�:���1���N_%��I/u
��'�L�����-ÐP�ZjA��5BH���j��D[�]��dx�s�3n�謣*�À
�@�1�U��nM�mA��'�wN0��dk˿�l.�gnE^�l��d�W|g�6����j�W^��¤/s(H�ѹ�Ls�j!�����w��F��VT�0��[������($=pF0����R�P�l�����k�C��Dŝz̦Vw����˜G�UV�3;
���bL^�A)/�K��g����G���C�����e`���PJ<�G�����bz����x^7Q��V����݁��y��C�!��4D��fGM�*۲PF2���L�r���:'�P����n�{��lV��A�
����!��$ە�@�$Zl���N�+3$��2�����.���߅ꥤO,�.| ķ�D
*	6-/��x���p�{ғ�]͊/��}<�DX\�y($#�O3�dy��~S�/�������w��qZ��#��U-/����Ш_Yp�t�56��품 &z4-�`�O��#�Xf�g͉;N�bV�6���I;V���6�zC�Set>ZBW�	�X���f����;��
xەY$'�d� %S	�f�2�J3���c���:{�o�s�5���.����np�dvA�n��s��el_q��+F"��ay�y h�^d��4]!׉$+�����G5������!Y�\���m��I!��%G��Wd�m��ga�U��+�fʁ\ٌ��Q�j5/�m��sp�D�)�I4����P�K�#ԗ����z��N3?7!�R���;�ƅ#8����(��	����1��0���-7yv����:CL��A���'g����	���h��5�<�YN$�{
o�º����LĬ�{s�-M��Y1*��2E�2H���TI�Ȓ@^D�JS����U��/��~o�$�#X^&Hx���I.����02�^�k�}R���vu�*|���bw��R�Œ���P�v�	�&�� C[�(
���fd������� �\�m%��f�����^ڃ�Ӭ�8<��4�or��{��/LS��x]
����;ͽ|/��s��p����KKRɢ�-jْS�y��d�YF�������XJMl�"q%�L�R��.N��p�;�N���r�{��`Rq�K.ø�*�. X�LI�����M ���l��\�M��5;2O�u�M��W���v�Q���E� �-�7a#.q�o�Sc�h���X����1ڗ����#��t�����N�wU�=���W��)vj\_��[E*���8 �T�^�wZ%������j�~f�)��`f�/	S�1J�n�������쯢/}��/I�5S
�'��i��el����LN��)�Ct�h5)���BC�?G���1<�%��H�c�|0�c��}iR���tT@.���2.�V"�`��eG���#W�4G��%`��$���&���{���Z⫱�qz=|̚9֓�L�g�`��(�s��icx? &x��=��3F�NX�0FS,��S�Ⱥ���D���=���]w�8@�K��(�^JJ�ȵ��S��IYd�����
�����{&�S������b`}��I�5�&,A�Tn@+j\�h�8�qM�NI�R�#�d��C���2.H���Ϻ��b+s��adFB���4���pq��f�F�2ݫw���.�fWw�ZOg����u֗7l�MK��ΰ���s6�a4Y�O���93l�6r���w�V���g� �QC��X����\�%�����ݶq�	�e��"���&�tH���o�q��}k�E�#y�[4h��F��!%v52w���Dd�όF 2��F�2U|6j�RSɗ�@�~iz|�S
����I���I�fڄ�堮��c�n����)e�`�۞Ϧ���Į�+7��:�΄�έ0P�q�o5kޚ]�F������8�j�ߐS$�-���Z�O�;�czrE��q.��1�T�!+p(���D�l`]	�st.��o3v�.т�'� �uu�c�M����U����1�˃싉���v�
O��a`P�TN�@r/f�"D���{�S�c���_���?m��S2��j��>C���V䗅���٬l&���A(jʩ�6Z
��)�4Dĵ�/���y̩���mP���OЪy}�%u�����X�����36F�� �6K[|���%��`�����'��S��F�W��Y8����_	�$�ׯ��k��I��B�o�� 3A���dW��(O�H�í9r�O�����>�1zX73���J���$��0�8����ƴ�m��lmU����xG�	��:"������I͇�IU*ď;��Bfb���N]�G��7�<��j|�� ͈*-��ma3~��qA� ��x?��㬚�A2��*Z�������Ӡ�uG�4]cDY(-�d����`�BK�mmn���	��[c%�����B��X������S� � �%df��Z�����xϩ�4Α՞�vf���۷p����u&���t�F���W�����Vv*p��{�w��䊡ԡ�5���rG0q%�F^b��?x���gwmt��ng-\C�EYY]�TO8"�¡����ZW9�vz0��S��y�)z7*T���
Qd���������(}����Ʒi�여M�&���{\�b�^�ئ-i��<�V4D�О@=���ˎ�L&���}�ɳo�P�z���Y���>q�<IY�~�h�X��YV>�]�)@񅰰6�ě��s��a�B�]����i��rV[�q{UzQ��Kl�ų߇��������$i�~������Ga��	��4���,np��O�W7�q�������i�!�����.[О�ڤ��D�%�/o��~VI�5�m~_E��(�m�7tC�o�;�q�V�c�n�v
[��i�![��Ғ9}�<c���'lQ�P��-ȁ�{ǿ�J��L�����K�	��-��{���Ց8B����;e�C�I�<�G�p�oHW@I��<���]V2U1:�ԓ/ނa/4D��{�����R\:v��. ���>E�r�<��R%e�)�b�51�0��Y�9_�x����r+�wH�**��z�ņH�+���m .�D2�ܻ�o���ǀ��m�1l$Q�@_Nv�wU�S���� ����86�r�UJ�[l7̋����K�����J�%,���v�r�dn�űOl�\V��/@��6U3���݋}��v/����?��荰Zr(|M��� �X|�$^��M�7[LL�+ϩ`>�T�N���~�~���G��R���ֆx8Т)䈽�-3��u(~R,�]��"n~C�߿FVJS����4�=��l?u��	�Ϭ8�q��56�%Uw�C�g\ ���R�x�#�5Wpڄ�Y���~S�a�S�y�Wv!�#�v3"�H���HJ�g��se$E�W�֍���~�X�a��DL���-��ՠW��E͏�3�o�-�焽\t[�m����pe��u �������Q��u{��0��n�#� �(n{%�1�	�?��=Y�=��P��I��v"4�8��emL<n�Z�rNW���� ��C�Jn�pe")�� C3,źQS�~OC�s�Gbz��.�1�q��}�(���H��)nb�����ı�QJ��|ک���L`�g�Ǝ�'�b���94���]bz����df�s�O����^)�ǩO��/���y8�����tI1���}��k7QOl�X�������0/�����~|ײ �h@�@K��q�xO8}�-> D��G��΃R\'���o0������>m'<��s���.(x�A�X�p����.���Y���]aR(�8�Q����|����L�dX����,gj��^E~GCڅ��{C��O�;�D����hu1X����<�A�`q	����ʏ�� %��U^^Q�V�c���U����q��Y�U�k.!� !���;]
����Q���>(Z�wgYA�X�cD�Q�T�jm 	�@w�+a��4I�Nm��U��S��Tk�d��ϰ��l�H�<)&�Px��y
�q �(V�������Uh���q�VGx���y�7�M�3h>��^�!�N�
ozG���.���ܓ��	���� ���bS���pR[�	�+���X�co�sA��ʕ	��Dآb�!@n�P�\�<&��6n�'�]�y�]�{��V?<���\{�����%��tU�h~�����B��s��F�x�n8Ѱ�e;A��'&�it���k�d��K$@�Y�{�:�������x [C��l����<R(������(��z��B�]�&�1+ݙ�~ث�KS	�`ؾ1�τ����M+���ݍ�E!���{A���#O�R��-�w1������s�\��ކ�L5��f�ij3(�/��ⲳ�0�5 �b���Jm8�cmf�E�vX�q�N��9JAU��=�\D���r���58��������lj�2�N:����w�Z��5�����h��3��D�sa3���(% "
w8�|S��u�N�R�13��(�ά{t7��l �fG�q�a_{7�[\#I!"9`X�1�{��5Tϒɤ�2v�K,݉/�̭���ID��pIY��s��Ҕ��
��Ѳ����_wl��bD|A�ұ�W�X;Rh�!�a��$���6#��S���ͦ@���N��W����j�ҙ��t:�<�ҿ�5��hcA���!0��c�^@�LS	c�Xȼ�s����u����'rQτd�	�>��#%w����d��U�����Y��`Hܷ���)�� �"� ��J��́aA�.���2"��}���\�AH֓֥�Z��ˇA�,Sa��QeL����(�#�uA5��\��� T�uHg����E2�<~�R<p5t�ˁ�"{o�\x3X��g"�������;����'Q�yp�jS��ײD��x�)w��Rȕ���_aL���7�e'X�@&WǑn�f��贺� ���'.{a>=�>51rل5?:�s��ȡd�y�`dx��`ty�k,T����f\;?6�"H;�;�PM��yG����u���(�%b�Bؽ@�a�Θ�S��0�O+��R�Ԥ��Go����}�A�ޒņ.X-E�Q�M)�'s+���H�Y���T@"�N-Ug�[�9B�7��s�"��5��Lr�C�롴T�x�cIh��5\�Wm���%���E�Mp����E9��@�^����'�������i�mz��_B3,�J�j���_ǤOAi�:���
G�{eP�����V��pJ�9o m9���)hC��iz}��e��-7~�v��j�L���+�&�f��KS���+�ٕo.dY�z1ץYt=ᩄ�*�C)V�����Џ1t6�ko�,"�[-�����Bq��
�����I_qڱ��sV�Ӥt�W/d��A�f�Q
��KZكH�q
�Li�g֏iW����2J07�x�}Hn���v�O|>;�|����c�Y뽠/c��S��.��3�2�H���)�^c�˵^���S����*H{^����t����3�
tp���
���3�YvȤZ��@�����^@��U����Ŗ�L�$��i8R���"��H�B�9UC��!ۻ�z���y�Zq)_����J)س��%0G6I�1.%�;�)�����C3�_d@s&<��wH�����1�W�%�#l�u��)X�R�,��ƾ�Ű��x&1�@�-�X,LSWg�r:�|6Ԅ�O�"{�~������Ӭ�Q���_�����=T�>u������ ੳ���Y*�v��ٯr�U'7:�pT�uʜ�_�g�J��j�|FV,�EMA���`:�q͌�J�R�*"MN��u�Đ�d��\����b�U��~�_�[A�oy/k �L������V���f�9NS���]����ūM�/b��l��]c�k��'��]?��"f⁅B8艍=*�R�Z��FR+�1�UZ\�V�d��C���InEvdZ=�ܨ��nl���7L1�a��^���)kN�ᇻ=*qc��۽������U+�,o�G+M�ڕ_�'�u	�L���x.��S���	�w��U�����
��6�d�*6��-7	_��a��#/�����@��֛���O��G�^k�E-�Z�(����S�B?�)�s{��2�ݻ��j��}��O��:����d��o��<�򐓝,'���������"W�Ϧ�/��s3*
�X��� �u���%rU�|���S���Fؘ�
���>q�/��35���A-���}�cu_&�Y���)����R�e���l�Ş�nP���49I;�F�١���$�<1|e�Ѻ[�X�e��#Z����RU��ƺBO��y@t�ry��
�w^�S�)'��)	��8�Ez��]��+��3�`$ډ���CF���G6Q�3�JՁ��$�����e���Cct������e�2��c��xD0��7��x�^2�9���._�4.��O�@l�kA�_��A��c�b�f�N1Q�[�b�{���/�v�2����_� wj�K�Z��¬�Ct�d��@f~�P�#7��D��$΀	�ȣK��3'��8�`w8�hc���F���3���NXsh0Wx2b�}��}�H(�x4��� xg?vl��F�V�H)=�K$0v {���t�����\%N�~�y�#���GoH���
�+�%U`d�7
�]Ddr�O����_�9C`�ɟg�wy��bYGжk4	@��&��g/�T8��Z�C_���4�*J+�nϨ�ۖ��}@u���5��5�0���S�8t���l�Gv5�����Rb^�K�� �oQ��a�*;�=���rM�
l ��(�4v���J�,�&5�� ���#��O��xFΆ�`TI�X����i�cH�s�k&6��/�я,��͕pp��4��ꈋ̰-9�<c�/8A�gW��2i@2��{QM�}��@4;�Z�ƲT��yr��f������-�C9;a�#�*�>5tM!������n-��W�b-�Y!���u;Ȥ�)�ƛz�A� *�swY�+��b�.rވ�1Q#��T �T"��f����]x[�d�x�L߈�~��0���}6��ڜ-������u�X�c��]��Ԑ�8�&�ݏ0��p���3?�.�楼���3����6���4s£��@5��O���S)	��QKQ��#�X}d*�`�>X)Q�9�S�D���*h��|�7f�6�md5�@YN,�.��ȅN�4��٠�/�m�iCK�����2�w��~��.;9��s{O}�ѵ8�C�Ѿ�V��
�:B|�r�v11��~h�X��?�>�=�V���.c[�iYWH��9�cPc/���!�ص���q�}��ø �{O����P �pA*�EN�(^�S��ĸN(j�8]F�&�"I��R��Ҥ�]^�Z5��ٸ�xLn����G?�h;),�P�����T���/S��B���sSZ�qf��-���W�R��&/��y��*P� F���bژ�ms:"�y4�AJM�'�#����VkdF�w�öwf,Ѯ@��i���Qd�T�ŗZ�6j�%��zy�Ѵ���E�_0��A��9v��%��2�#���k��5l�o�@-��t�P�S6�Ĩ) ;e��p9*,�z�H�H���r�9�:?��!�5h�@��F8� _ !�lz`���
*z��f�2��g_�ц_lP� P�f��,"����l vX��!w0r���-�����P��׻w�A�$���p���(�fIH�L�.��bD�֡\zj1��L���{O�2c�
�ka!�;����+ͩ >�����Q�g�>ϓQ��'/�E �?��f�s�?��d*�G�ʆ��o�aGF�p��1$��T�^�5cHt��m&בuN���'�S�j���]�d	��Ќ �`�KO��A��&��O�`�/�^կ�?W
w˄���'�{�������[3�ư����e�F$e�2��Է�@��(� ���#D)��k�=%�/��
6$ogw�ZQ�O��< d�
�HmS$��!�f��<�˫qj�\g��[�z#�@�3?�3^]�L�����V�y1yz3�P
q�3e�X���qc�{�;;�C����|W��,��#���X��^4�Ä�R͉"M���x�����jE�]�0����8'�?M��,�czz<Ļc�W@� r�Wʓ`a���]�bU�% �UP(?@�7�E(۔�m}�/u3*QfX*�ta^:ѠpQ�3��_�cbQ�w̎A�����5����%75����\�}�M4`��L����)�Q'�ԟ�8P���`lJ��J���S۾X�.M�܍Ӏ$|s6�m��[U��Y%��r
l�;����k]U X&��7Ĝ�թd�#���$F��䪣6<,�=��N�-����j��u� ���]����C��{*���Kl�~e��U�p��E�n������<K�r��Æ*����i|u��h�s�
����d)0�X�
�IS����\"���M����#0ztw/�NF���F���FX���}��C��l/C�/�sYbI�>�W%y�1��"	�p�og����iҵu��'z��X}�4u��&Q��b$#ԣ�uu����wh7�p|�'I�~�D�w�k.�������s�z
��dYwAJ{籹������Xv८b�Be��Bɶ H�e��p��e�k�ۢ�8Ω����)���ɡp0f�v ��#��${r�������}�V kخa��>��ۤV�𫐖�4��`���'���#�j[�m���ί˖ן12�*�n�翣+E{��Qy�Ŭ�-���������ZH�R���vZ.��(a"9YjK%;/�Ql���O`)cu�ħb,���R�����J�.DT�Cw$�2 �ʌ������Կ����He����M$�1J�kk/�����	R��[A)�]�MPF$� 
�� ��5䨫T��[B���6�`M��:�J�XaGs��{���V<#�80�M� �s�C;	D�N{Bϙ������]���Z�.(h�gPLa���=�o�V)^8��˭�˒@2mre0$@��J�5�6>���t.��u$)��{�A;k|�dx��	¤ij�������ù#���O���̛�2���&yWǕ����ӺXٜ�������P>�h-r:Jm�1��p:�����w:v�2�،���~�c��v�uJ����L�0D-ޗSI�f�8�(�}���Qڦ^a'��G�:�5;�5�/N�:]����K�q�A���˸���z'��E4�B�
J嶔��qŘ���9��/�Ԏ��O$?V���:xJ4����j�Ds�Ә:;$Z�N�g��5+M	�\��J��U�n��H�[���D`�+U>��{�Q��8��h���B��
�a<�p�A���*s����������C1J�.�q��=6skf�ع<�;�Sh��G�3=�F��v� ��n�p��?2�����ȨO!
j�T9��������?gt��N.k�RJҪ�I�>���� `U �H�L����T���' �S�r��k?Ôw���.��n��z5�Ak�ﮭ)o��f�o-c<[��ĸ�N`.�~���ڨ�a���>��}qݙX6��j�1ՙ(��*�s����ʄ���{��D��h]z$C��#�Jd��<��p��5�w��s�AWJ���$�����;�)w$�ѷE�ӡ��p�'�~$w���I�$�*H]��,|8�壽t��ݬ�m�̪���m�O䎪���l�/m��lF�Od�}��dIc���hA�ӽ5�|����\�>E|@G��5�Ω	H
���S���a�هR��1;���x.�+���d��#�G�����v���+�$��x"��Đ/q�`T����O
uM�'�@���q���[W(�����}�4�0^Z�1�cWT��(�BD1��}���7W����c��j5����w���m�*4ϵ���)��P)�.�:�ꒉ���U�Bm]?N߭�_�B�����ş�N����zv� �6*$�-5����m������>jI�A�2�ZI*�3g�Ɵ��(��K���!���u��tҧН:2a�\������Xq�?���܀��%�&�b)�h@�=�V@��NRJ�?xY������3$�A��Ȫni{�������˶�!E���l2^�HSk�R��V���V��(�q�X!@�V�%L�L9S�/HKRo�o7F}FgB[�q�g�e�ᴒ��P�.`��l�a�����I^���>�K0s�Dm_��w��l��xm���i����5��:'a�K���v�o��0��7o��sE2^Xw���Z�,9����c�r�L��o�<#<������Y6c���J1��e��,�Z���z	�Ҹ�RS�2G��҃~z��	�f�%E���3�M���-�Y��-�!x�Jg�0���?� �O��L6���Op�s�y��i��]g���6\)�cș8}����=P����Stq���'j��TE�zt�P5	�'��k>��@�K8*E��U"'ظX�v��d{@�)qr�;��\C_�Y�x�a?M��э�;�7L���p.L� �$�;�#ڲC{�e��������J���Mz��?�|�� ±%q�u�����������Z�R�������$M�����8��3�:�k-L�(����I �GT@ŝ�?�~�l)�N�"���b�m��vƥ]ǧ����ti�3�Ŝ���D���?Ȣ2$	�G[;O��/Gd^���ƈ"\��\'����(�����j[o:}HU��b��� �ԍ%śR��S�������P���*�I�ׂy�0o,�"x��&=<��(�	�{1�[�tUF�I���]"��$���i�&D��H���sD2��/\�ԤwnK�{����
U��A?�4�I(�h��TL��t���Ӭ�8֎s�º�ϳ�>W���W� �������~�W�i�VD���$��@�;�;��wZ�ks��̖�}� ����:�{A�}'�f~���rk�"�Z�$��P��h��%�j�h�`٣�I��� ;m $г��{A�&B��A�(L?.��a��&�vCr;ccE�oI���7>��ل�A�o��<�{��L�������J����qy�xm�����w���X{�kώn杢������O�B��Wc�-�r?a��|����`7'�q�������C�o���j�!s2�G��
����+��c�p�M���XC�i�=	�y�+����b���?p%pR7�?�f������	z�]b4�>
LTLn�=i~�]֕_At2)������_������m�O�Cy��b�����1k�x¢_��xEw�k��-�h�Zc�%��{,���}����K�`�)�#�����K"�@TO��u}H�Hui�l�{ڂ�3V5��_v��v+�O@�� ��̴¯���};z����J���A7��b�fU�����- �ñ�@���P�7q]D�������	���U��*��]�L˺���6�<��c�p�3ѭ�	O8�k���&��ڜ`�?9@7Hnmv*�<��#��^����Z��s�r�����b�٘Du�"b:zS�G��%���o�[� D3Ӷ�A6�,N�3��&}�i���(牻6��Z���w�Q|h��z����V�WK��!Yy�1�����8�蝨���b�{}��Oi{��WXb�o4rKJt�Z�}��~^�n����3dn��@O�4�eHe�'�=�H���q�δ2%��k{,�[�N�M%YH&T�D3�J��Y�o�1l�n�h��`ң]��NT�G�<����؜�9��҆g�1��h .�T͸,U �O���#ઞ_x)����ad~V���^b�`���e����rH@��/8j).r_׎Z����S~>�D��a�$�+ѯa-o�b9z��j��4_��V �W�7�W$����љ�r�����;祜u�Տ��QN����R�YL�;#0�����Ҁ�!̨�F�؍�D%�N��e/]�x4b����Rn�O�E�i��AԞ�!I���k�6�S��-ޡ��X��W?X$�$vA�Ah�>.�Ih�
�T����7F�K�,�䴩�C����ʘ|L�uZ�[�"�q�E��l�&ؒD��Z/7iD�����>�xL�t�*W:ń��uF�)Ϊ!��̮ѢҞ|%��,���S�|i�y+�6!��a�%�q��J~�����m����Ñ}����6@��=��}�(n�!���4na�RZ��^�B~7�p��׷�y�j%{�6	���A�ɭPu�t�6��]�`�V19+{�R�v'`$���d�l��_E���Y�8�.|�5j�;��X(q]��Ta�h	G��Ѱ�"վ��N�%�����mW4Q��s����M��P�Э���!A�}��Iz�NzF��hu咅L�K���ɠ�~���#F_���A��ź�f�h땱,�AǴe�����a8b1�(�HH+2���|�y!��r���a����vfLu�q:}��i�azp��N�@�xn�Lˇ��D2���|뼯#���H��Q���W�~S뫋~a�rW'xN=����NkP=����_�|n-,F���X S�/��?��Jy��k�͏@�n��ҹ�a�y�l�M��g��kظo�N����L�[p7[VN_����v)W�Mc��nZ��ۑ��xn��3�W���D+�1���5�?���&��Z�EBT�d�^K5�'@vs���	��zmA�nZ�VfQ��wn���o�c"�TJ����C��B��,�w_��g��j,
}�Ч�y�lA0ͭ��z{�w+�XN��B�-�!���vb�}��oi�g4��3"m�7��I2n�v����zW`-��ɐ~cg[Y�vC��u�S�<WCI'�^ƚ������T�WÈ І��t���w��������kM����&�S��Is��"'C��� JWi�!�o7lb�hnf`����碡��#��g��s�>�J:<�N���h��L�jL�<��˷D�|Uה��-0FK(�B,Lv��OҌ�k��w�g�ZGߪ�Y�
�[�p� �Je<�5�0����6i^��Bj��>�*%}��+|��7�lc�,�f-�,w>���g!`"?οxW�R��ȹ#�e� �¹H΍��~=�H۽w�~kX>����n��!�/�(:$^|��6
'����6��,�����7S�-ŏ	8���ymL��k�2���m�blE?�2P�5B�l�]�r���]���s��%�2�4��8ۘ�����6��uϳU(�vEq.�K_�`bT�ؿ@W8�ǈy"�p+�(�7N�tS@�խ�~����0�B߹������Z���g7�l!n�����N0
� ���X���=ng��L��F-N���+Y���|}��,�%���2Bp��|���l�����&l7�)��Sf�Xl�ؾI�d���n.!}
��)��(z 8�3� ���02.�j=u�p�"��,��sc⸑+���M�y)�/��ӊ&��RbԳpX�� ��}�{w�HL���]� �� ��*���\F�����qܖE��H�DMQ^������O���1ɸ���xq�?�,FZR����O��B�z&�T�wT��&��Z5�`0$ڶ4�T�ޕ���D��<)ф�Ϸf��4B=��mD`�?c�6?7���	ј
��g�l��{ ��zi��f˓:x"�/����R��k���@��Pa/wj�s���($e�xэ�^�C�?�!��e�J���G�N��qLp�(�q��2~��F��>��`��Ǆe}"�ŋ�ˌ(��N��>ڗM�C�>VD�H0Z߫uy�'s��{1"Ƒt��^W-Sef�$���]:�}�vtq3��BL UEH[�J��Ĳ�!�����Zwzk�l(���KLh;QH��ʠ����_M)��g�t�m�`��y���)����f�ֶK�D6U~�%5�� ��=xE#�C���M]g)�h��z�O=���b.0"�s�NtDkv��Ex�^~�D�#�Wq�n��c̰I��C��a���RҐ��MF�/So�5O� �0 �F��	��紐��YH1�x��<�)*��s����<�l諘�Q����e͹��ᮠ�����{hlnuM�{�4IKr���<A��Ew���
\nw�O��k<t���ń^A�
�'�fD���.�[ۅ�hZ�O��ă42qMmy?��Rb=<�ly�G�Y����}#rMŝ��.Ē��:/{am=�e	�r�`�&��}V���r!s{9���d\"	-��<<��-
|eh����|*'J��������=_5�rv�-j5Id�l����7���j��SK��C�J�g����Ec��3�}���jCA��x"G��Ϯ��v�U�18��	N��ǲ�l��nt9�ujS�� S͓�*z���+^��u���q[�k"ڂ?���˯�5��@쪨X������ .X�H�L^��c�pVhզBįY�	kHs�.�b&'���v�6����s�rU���3X� �i��S��r����}hI�^����(sE��1�ӦAc���u����3I�����L�q������T��\,�Xd�3�A*X�HY�����E_G�`G�H�w!w��nb�_�򊘒?����-��H"]���-h�!�O/��mO��l�#v\(�D�8mS0Q����As,U\�;��ġ8�M՚Y �X���i6Mi�[K�'�(�e����O�ܛ^��6k+~p<�z���Bw�t|���I{��'�e�ե�����,$�G�'P�*)K���G� ���}&(������d��z�\�0��k�P�c(9��y�Ο��\�Ī�k'h�^�ܼ FL�|��C��0CQ���f0ڀ�*�9�bS��]&���݂�t�D6J'��h��u4�]�1��9�jd��,d� ��ZZ݉��g�]��m���"S�1;��"��h�X�kU���4�� ?�qv�g}���J�wī�?@��Sd� �ގtV����*���0�Q'8j�C��Ӧ��	������o��*�g����)29B�����X�3���5�ֳ6���Ի��:"֯<p(q�#4�2��D|�t�f��X[���y�93֙���
���S��c��:�/K�Rc;�U�g��?,�D����M �+�T<`��]$:r��`��m3���gp��3��:0�m[�������)�fp�Н�x[m[�Yڥ�cL���k\V�������@��[O�Fc�!���q*�?�U@��-s���3O���Q`���6�״+����a8fPP?�:�;��zo*�'_Ȥ��S�����p����|�0�:���?$A�S>��Xq\ߴp�m�,�7J�̊^Ŵ<��lN$���n;�!�������j0vK�4a�yϔ˩X�ɂS��CL� ��-([�X�aN�VM���E&�SK���3�i~'��cKSy���Qӧ���oT}��~.'�3���p6a�]`������?Ē!�w m�4\y@k1G�F���AL���|<�Bu}B��Ѻr����&�V��:W)��<c>N�|��ٽ��B�9�_��@�޹k�:���#�� ��aU�����>߬�F&�!�h���ny/�`�[��KM�A�x JQ!��L8[�����������/,�w	�9n���(�~��~�~�o��,%��?��m�w�^�����4�dz�5����ST~J/4<��2�P����x��39���CZ��	J�1�.��le�/����k�]�i���zY�|�zݒ"E�Z������P��0G��#��=æ���X��W�ͻ��WYwY|���Tʜ��oD2���+d�qd�!p�G���ai?��"����z����b�j q�]]��^~�[6΂��6ᠭ�G6�����Y��yY�e̛��q]�W�]!�6+V˂���ď2dJ�{�����6���?� y�4����S4� ֹ�ɑ%D�u5�Zg��$>1 _�S1��_BBۨt�`Ր��㛮�hN\q+���&��W��j��t�{�%���pAs�y|8�@�)ו>_�+�C���W�[��䔯�8�=�����8e�)�
��n�dI}��>��C��L(N
��5��#�X�ο��G��jR�f�(�E�6	�ΑM�Q�?�]�T Z�����Z��ݛ��RD�ɘ��i���M�#���o����e+K��E-;��9Ro
����Ԕ�������� 3��.H`���s�lLX3>O:	{�}]���=o,la������̻H��6x56��ܺA5ٷ�"��+*��"n)`
�N�ةvJ꜎=��&o9N�Juc�;o�;i��\�"(�������On^~i��' ����w�[[�n��e�u>�Ǉ���5�i�_pg>�P�F�w#	B��Y��2˪�ɆږbLt��1��d������|3���[o�}Z�h9B�rի+rd��D;�M4)�{%5f6~fd�	֡�G�?M(����;9b����g���4�a�u�:Pn;����>���W�Ș�W�Pp!�V>Ws����	�ܳ�mk��,e�Bϊ3�)�J�7�Oip8$U9����t�!���vg�Kl����C�
�w�Ͽ�%�:���,v��7k+���ys��m�s ��5���12���Ϝ��O @�"'}I�ھI���2��R7������?���mY�!/�GB	��?Y3&�N��X���N٫`B��!�x{����"?:���Tӑ�N�[�w���[��1 ,��|� �v��+K&�{��:4��ۓ�g}m���H�j���d)��Ħ�� S�~)��cj*���C孅ilc��?1�/:^��4ϡ=��z���RK��܏f�&�_��ĸ�S�����$F�H'���y|�+7�V(�[G��}ny��_��jm?9��ظ���m�UnF����+���E������"�����y9�����ϊc*xh=��J� >a�?4
W�k�+٨!�G)*�4�
��"�KoՊ{�G�^;{`��(ui�b��L��W^E�9��{�y��ξQ���f4e���՞|,1'e4�Ǖo�h��~$k�׆�E�d�G�Zڬ' :b^K�`²�M�$����y9o٣��wk�|4��d������x/aT���;C-��[����R r�/���]`ן����>pR�X�X-I�����ȇ���=�Rz|z����J����>�\�מ��Q��	O2��C��qX�s���ƙM L���ѰOcq-_VW�<"�2*�	��M���8�y���tr�s�eD1��jF�ћ^_#����Ҟ�Vw� ;c�bb
M�os�>�ȃX�}�"�f��1p�=M}-��*w���FJ��B�G�n�_`S��޿�!�����@��d"JhX�\��u%�C]��u�X��Y;��W6��� ��!R�dٻh�)�z��UM�((-�}��������^��D"��A�ێqS�\e���=�뫦]6����(�#��w4>\	�@D�b"0utC%�|�r�2q����	ݕ���>�W'񎠞��;���u��/�?�d�	rzP��%��l<A	��V�vw�� fϹ3�B�x�D�>�L;;��p�te��m��B�Մ�GJ�JN:�r<����JQ3PZ[[���L����Q1�f�%�"#m8�y4�@�Dg�(,0 .�K4�~�����6�[*Y�J�S>Z4�m��?�K>�I����D����]�d�eU}�<=�x��@b��Ip�/���Hu����o�Yo��	&�e��˔�L>r� �����Y
� ��g����g�@u�#_竡kÕY����J(��$t\���v\ўb��L�;U�Q q�x���_�.��,5��*��B�eO_G�<�^l���n���Eޣ:G���\��6�Fq}��)<2�P�+B��	S�B?�C�>< �&�3�;��A:���m�D��$M+�1�R�Xo8�clB����lU�V$9�"��}�.��  ��ʽ��k#|?\�+z�{BK��Mг�]���Y[�nݜXao��n���=t�Xl�H�R�U�9wt#1|_�+���X8�L*��y/��j��E�Ƹ�qkb\�my&#����Mry*L%�.�3� �#����;�~�������� ��#(d�ʞ\���s���T}C�`(j2���UMf���(��l���S�#���4������˺��C��G$�~�����v>�9g�1�� Y'yW�PE�բ��!�S}w�\S#Y e��!����$�`����R��y	C�j�d�0�{<�;�;%��}4�1���ɸ�%pp+�t]�����q����e�[���I�ETsԮ̓������UպƬz�"8���:p^�$U�e���v-��:%]�Q��IyiMH�9�>��/����m	�Ծ�_P�w���E����I�$��"�P��?`�C��uFa�gː�E>)x�"�0@uE��c�%�������W��X� ��2^���|�p"&���:)�F���*��ȴ�,;H�M�c���[ܲ��O�[�R=.8�8c�LK����w����+��%���ZI�Lc?�Ǔ�i�Ѡ@A��cO�M����`)ܿ�X:W �|0�_�H����?O��dc��rmk����X%-t�P�ˢ:�-���+��bC���?��y���FW��d�+��j�a��.����쐃J�+Y���MW�˕�XG�!"rxl���zC���ɞ=�y3�c�B�r���}�ޒ�M3�2�]�Pp��q���@ ��T�R�23Si]�K�{�+h�v��\�� k���Ԕ7�V	�&�mq�*�AY���T�?��=46��4�:S����+��vC����"����'E�y�n ҧ�>&���2����㔣�Bk��Gݳ<��s58:�f-��2m���}��S=�#tC����?�E>��n�$�,]1�:�=�C#��x
�ό���㏄�v�0a�d��)Gs��aaI�I����`(�9N�|�@(��yO��tb|�TPAA������Z?G�뵣*�k�?e�C��D�)pj�.�m�9��f���Gi!V�7�D�Д��3��KtG�f}����+ӧ���X
h㌀��T�/��o���a����sd�=v�4WF#}�*3Tɢ����VV�	��/��$��	��F~�d�{��;�bXo��,�G�:�C�R�bi�Ţ	^� �;a���v!8��t��n�B�Fv��Ck�hZQ�FF��Q�_'���x�{���+��Їs��{#w�� �(�Q7�l�%���(&�o������0!�$Z��G���i���`�RB����yhU���,��#wi�F6$B��R��c��������_��auIu�,;|y�+/տ��90���L2� �PS�j�y�u��[�m1���Vq!��	�1h�#d4�n�{��q�D�@A�{C�[.?��yT��G �B�x`�ܾ�e��er�ŗh�3�ߩS��v�8���HzS����5oy[�C�3Jn�Jd��u�赦K���i����7��� ����ۋ#���uj�j'b�a�Q� �"����x=<)�de��"�i{!]��\�Y�t�ր�sںf�-7�����Ɉ��~V����	Uw�0Ѿ��y�~</�>�� �����������Fv��^��T6�W���S�EM9�g�8�ƃ8$���	�z朽���'����<W�kg�]�`���6}�[����Ea�u!ُ���o���x0�E!��J�[:`D��o?��^����8�n�' �a�+hq�B�0
���$��d��o>�� ��>ڨ),0>RL����J=I컻�������L0�\��M����֏����&e>�k�����FP>r*���;�t�U�V�&�2l�2=v߬�l�2@ױ	���e�P���c��L#�CO�%5���p#Nt	"�|��,d�3:?��8k� ��Q־@Z/�O	B��k��Ŵޜt���6���ۜ��#H��n��u7.v-��>�v	�M>Z��1#�X&g�	V�� ��Yz��5Um�����;����i��X��T��L�f:� ��Z�N	(+v%:�{?� *���s����\ ˣs���n��5���[��(X����һ�� �Rz�NzF���=䴞�[��*� �t-2��v �Z��dZN�߱��<��9��
�FB�����Ce�`W���$�J���f+��e�\����ae�*֙t��ޚ��Nu��;U�L�צڄN��K��a��crM�#����(±��5W$��qwT �q��+V��\ԓv��	�&�����|B���Jmr��	���fu7�z�Y�^��yl��Pޕ7�7�B>6�_�n1
���2�����©����6T��6+�;��jb)�i�BY�.`d���^b���/I!t��MY3�/	َ�EJ]���1�L�.0����Fed?���+�Ft�[aL�-�<�#k��NjlWO.(�<��/���1��IT�D�p�,x�t�q��B����Wܡ���R.-��2��}o<��P�vrU�����W���\	妑U�1ý���t�t� �U��~A��m9�݄t;S�a�f!��u��u��~By�5�1���x�@��;Vx�@R�
w;E�Wa>��VLJ��T�jd���{�Ə)� yk�3�E0�Ƙ�(y������rB\ ��48y�4��mo�*m��0��)���a�e/�����o�v��V-选=�`Ǯ�TUH�d���g� &qN����h<uh�C�����g��!\��+!�
oɵ��<slz��@�O�4��}��/�[�ǁܓ*�C8�:�L��B)�oQm�;U�s��U֥��>`�uD?鍊��,��~Fna^I�Na�����=�ƭ��ᄭY[S�p�y�Y�j�a�� �lcΎ?'��Kc'F�
�L�@�J�T�k��ڈF[Ju��5Jϥ���x�X���O$I�F��d
G2�|Y0I�CWʥ,al4xo��J�)�� �)�Z��g%�2=��h�G�3�`�c� ��3�SQѯǡa���[�Q��Qa��m	eK�-�}�Z�$l/A+Vb�9N���yb�7����%[åZ!]�d�6(Z���ZB�5U�rÈ��O�ǃ��3�g����s��vH�4ʏ�Uy�~�;���&NF9!R�t�kS�&�ri&:D�称�Q�h�˕<�`S�e��4�c7�.Z�N�a��|z��|$�a�yY~B����C�PZ���0^de� +�%�ݪ�B��"+Ee�n���i�fu�� �g��4$�!w��`a��aH�Gc����yrj_��>��ej��Uk9kc�/Z�F���l���M<�UYbS�¸�@��wr������ہ%�����~��E���g�ht��16���#�ls۔I�2:\�\�=�R�Y��7��K��;�q*FA�T	"��{:���|TTe�P���[^�L�L�a�P��x�p�Gx�O����rv��Es^9(W̅�}�a���3���o�k��2�X9��%��J\u�q�B|��HX%j�8+"8R�*m>!����:���6@P0`r���
�����b�R� �7�Q0���0Y�P��A �9Ҍ�]]���2�����ɥp���{,�0�P���LKp7�w�n%����.�y�3&�?��	+$>�P4
8p��� u���66.4�����z�Gv}�ѫ<�S3Uj�'
���Id���U��@�����W[Ɛ5ʎ4�h�<�O�y�!qGG�#!fQ���`���'��Ig#3��� ��}Z~�����G�
V`�5f���c�E�J�����.Iђ�=�"��dB!�3�B�Dkז3ޞ�f�I6�8k�]K@Nm>���L�����h�EK[o���r_n��C|�Ȼ�aBp	o�]n\ ������^x�+d�;1P�}�x�� ��ߌ�zg��;o�����Ad��k@��._�~(v<�x̴8�s�/+:rCFv��� ʫ������D��>V�;bID���1���:{Ұ�$K
�`�/��
Y�+@g��_$�<�ZYʾP��<R=w�=�8����'l�7`�E�j̨C���?��@�Zk�<��i�Sʰ%9M��R�&!r�L��*Y�|%q0�^�4s����q_�����G?寡9�>t?B#�޸>��~��-�Ʋn5�Ə! ��"�&y�<�x�/��I�Yx/�@<��K䲷�]�bН�r�O�mɏ�қPi�w4�r� 4�N|8���9Tݰ	�tI���0�t�|��b>���-�����ђ�B��b�^T��{n���0��?B�Kn�Dt�4s��9 ��柳�w�K��L��F�D��6ӻ���ش�Z�*�&Ko���2%��u�,&���L��G�E��	<,I?-i�U�{�	ۀ4<��ɳm2j1݂�D���=М��/P9��a����e��5��w/�-I�+�#�R4CGЂ���z��	�ľ�6�
v�_�~+f.=�ǫ���8��_/����_��]M�~��)���S��K���b�P]�@y�nY����G���Eӟ��7��\���ZG0w��W'k�V�ZD<�su�ϯ�m�[(�i���n��QC��M1�\ͻ�Z��s�N'����N��]���� ��齋�L�a��dK� �hʋ��!B�y���q�59²�N�;DW�!�.U��NqL:�̹?l'��iׁb����P�W�r�7�a.�#6(�~z*�)��V睼�{=ZO��M<�#*�O_ڄ=��	�&��34_���Dy���Nv�q�����B�Z���C�s4s��g�ۏ��K�<#1���J;���&B�T۹ri�܀҅��I<�%Ս�����SK��d�O���ǴA��L~�;7Y�|�0=$�Q��F����_���~gsU���ي�>=�:�	���r*SF�Q�̾묟��^�
h��,��M�#��/�Ѹ�X'2�S�Bb�E6�ru�0%7���/�C��Rxr��F 쐌�gc�
1�C]4���PhM@���T QlE�=�5pG4��:Å��_\+�Ou��'J���
�|�@%
7:�R"��
x.�/�'��$���a�h�Խ�|��LU�Tj�Z?�f5fg�9+�+����Ў�9R�%.h��=嘼q8���_`�B��6�圅�������݄����\:_e����R�^\}u�ܲW���?�9GmCM�
��4%�J�75Z�=�(��c�h���)�R9���/)����[��Y��@�I;�b���:�=}�/����� S/ژ�S6X$����
� �R+ڞ`)c�	�߷������|>�K{c�ps��XrG�f#��pۦ*}ȫ�E�so.x�"F���~Y�WLr&/߯%*g��0����}i�bR�m����Gn[lu���n��� �Zl�?�IS�X���8쿙�{@�Il��Ja1�fEs~�M�l��\��\B	&N!Ón(X�m�W/��彻���Dm������-�k�s 2���q ����*��ܶmuѤ�V�؃`������[mݫmm-o��H�c,�p�M�S|����� �7R&��54&�lg�!����ﳺy4����Q%���r�ך�' `����ċ�B�5]�̛`>-��������V��ѵ5.p.�SΘθ�ȅ|*u�
Yg����e�ffO,͚���z�
~x�Ȓ��֦�W\��Z�>����G�,�*yi�	�,r�h�5��ȓ�"6�s��#(����6B�����P���u�3��
_��UN+w��ڝ5�9%S�!�nXn��t#��w� �=�	��2�w��#sݜ
�5���h�.cǓB֬��s"c�e��wq+�ES��V��4�k髴�q@�w�f&�(��7	��M )67�?T��c�v8x�rԑ/�k�l|�O�n_V� yR�͹�#�8�Y���j#ܖ�Eq�b�PIERx8��3��H_��¢/?�lC��_h���=V�.y�q��V~�@][S�Y*�a��h�CK��쭨�����Τ�&�L� nՂ[uضO��+y��t���0�@z.�R��3~͙K�Ü��0�jR/-�@���+��#�~��gd��$�bY����z�\���h ��O|�By�s��9P���Z�ؑ������t����9�а�y��Ұ�����O<��H���<i:_i{����o۴��Pg��i��x�!�t�zKrfg��شk�
b8ʤ��3���$+�مgNH�oy\��r�T�[�g}3��br�_bAr��1L�������l��]v:~_ДNÞ����������ˊ��JC�/�]�z�����J�5b�}ڥwI���My�<ߚG."b�B>ƃR�:J�j�ǅ"<��29�����̜=��Q,<�:+��F&pd�jWtFog��j�MV�|&U艛;�������_HQJ���V�����Y6�k�T��ُ�>��C�{B�]��K�EH#���姂	:J�p�������3^r�
�~hЕ_F'A$)���p�{e��cF��B��E��*�8��c��5|�d���ZQ��E?��}����m��?b�'�i�Cz�Ϙ���_��M��&
��wX�UUQܾ1_�����Vh������������o��7��ׅ{P�z�x��߇�t��/.���2��`ɍC�^6�o���R+������	�tw�Љ-P�#�W^3|Rm�|u�=z��3o�"�����݂�7f�4h>��RP�c��|�Y�Hظ'��J!��f9k�j;Eܖ<�-nE�fܥ2��Y������?r���h��:|i�n�"b��RX��u~,(��Zp���
����}�(����YF{(U��-{�n��ˮ��A�"��oSϔp�jyp���J�2Q=��j�tH����k}XM�AX��A���S�D}�w�p���rw%���ՀXPAje�+[7:�)e�>z��ȟ�4�d��-�ٵ��E]$�P�-�~`y`���u��l�LP*嚑��8_��[�r-N���UF�[�������m�=�hOV�RPB����Ӛ�(^��ȭ�<�m=�+��˰ES�p�O�0�\��'��8�R�|���Ѩf
$��pf�I#Z~w�{��#���I��:L�X�~�1�"�R���<�q����~k���d�P��s)���a^�'����~�dJ��:`����@�͖�k򱀺�w\��F�E��ۣ�֨U��6����
�(a�X:�����#�c�dXk�B	���{.s縦��k���i�^��TE����k7���.-]YI#NH)���
IuS(�ۂ��.��,Z��Ì��5�h��3�23Ga�G���tlYw�҈�� �w����Mx�5��;�⎙���ĝ )w�E�7s�d�c�|"�
!��'��=o���}|(��Ukp��۾��ڰ݆e$�1ch���6\Lš�
g�s<��h��?�[��c^Uu�%�Ђ �[��B5��m���`'��[r�0�?zV���7�؋�"o%�M8��Az��σ�F#~�t5��G��/ģ	��sm5x��l���]�%s#(*�{�VX1���k>4��5�?���Ӈ�c�=�S��t�`����BZcg�O��)_�*�gev���iT�g�pq��i�~1��M�s��y���J�d`�3d���-�Rh�sǺʡ���C����C�q˃���F�O!0���'S�"8a�~9����d�*��E�+\��+)�@����V(����+���Aܝ��x��NAD6(2����s���~�!D��>�]@� Qr�U�PX�p��v�7ێ����
ڧ�m�} �MO�Y���Su����k�7�������K�A�+��*^J�P%P����1�~�|G�P��&%q�G/����˒�U`�����D���p�jo��+a�&k�� b�/���n���� �ޱ'[O���;<�l>�*�h]�J�=�j�[`����Z�,�����x䠜o�'>M��Z88�-�$4	(],�E՞�ESy�th�!ޮ=��#�~]���𩰏{u����;�@m�p�N�A)/��$��?ޤG��Ҡ�"|i����rHN�L�*m�D�e��sI�Đ���A���m��r���8�?�~�5Θ����c�f��.o��.7�A�eߩ2C;)Z���mݼ%� ,��)���U��*�s�VK�Z��ء��H�J�=��3�x�i5�W��{ {qpۘ&�Kt&�U�4x�k��W5�� ���5�ʑҀ�b�B%?Љ@K�r�1��[�F�����E�n G����T��Pj���w*p	Z�i,7���qlTC��I�h��elUw�����RKN�#�kG����Y!�%~J�z����G�wƒ;oL�Ц����$AlX�%����{��oj��*[���Q]������o2Hz`r����X��1Y5�[�!O>U�H�,�u&�E�}v�k5��E�7����Su��A�p,����_g��N0	w|�p���� �a�r���P����5��鵙��@U�����oζ�:9a6kp?�`~���䎕3�PS�	2��VS\LR\�{$�U�F��]����+�;-����'�?�f!zR�֥4O_2��p����%�.o�g?�9�.�}[�� }�F 3g�������x�F���/�K\%Va�����('���?�V�T�|Nͱ%�$���D�Dـo�
�~�4���ZЄ���l��E�0[eu~� ���a `eR�w������c̟K����yͅ�g{�]�K�-�M�ÁGf�Z�H���#���r���}|(���|*��7�����M�U����As�\�88�f��ie���5D5�}sq�$���n^�RCyپ�Q��a�U5��^}Q��i���}�uƟ�8:� �]���fz)�V)�n{*{]yM�[$��> ���F���Ђ�֯5����&�Em���-]Ӡ8��ﾤ��_R��'��Ǫ���`揞����6M�ïu$���&&�2U�����ًb¬����[ȃ.�����}�^޳,p<v�qj�D!��mP��׏| s=N����	�j�S���u�'!�@�#2��8/�M0���R)������l��!��%8�VO��dSj���H��(-�c�%�yR�QXDD�|a�n�>}S�|GT���~����2,�zH+wV�0���un4⯸�,���I�M��,�n��l'��(�HΤv�2�T\�� �٘�Qq_�"������Sn܍�	�R���Ɗ1M��nl8�M��D_�o��|.����>����(*�QАf[k��a�.K�����MkK����o+��{�cr�o#�{#?+$s�s��X��a%q�bb�K�k)!��]����q5�\��ہ�����<�9)b� ��q`�C@Z�_�'J�CV�j�_%�#��0,�@_$�B������S��v�maRc�WxI2�F�l�<ñF����{��e��j��m��ɘ&���Q79 <����|h0���Ӥ�#���L��:��>���Pۓ����:�T1"�����*�m�}�(a�Ewh.�V�\�Cj�٨+�7���Q��/�M�N{�6��n���/S:M�b!M��W�� ����2�I����&#%噂d���A8y���-Sx�~���� ����/�G+�2?�o^�SC�G$������D	W-�<R���H�xyK69��G�^2ng�)�_3���|T�������faĹ�W���<㇪�~�J�&�_�0�Ϊ!_=�P�9��_�bv�4샰R���*��=��_�Y �c�2Wi�B�G���Nyo V`�-\�����~�tG$R~4�Q߹U�wܣ��� [	�:E)["�����T���'�����\=�D; �%�r�v������	�����tY��+�a!�G������P� �@���W�~k�]�ޫ�v7/f�C�(�<�"��*w��o/��А��� t�S;fi�,�'��j�yR�J���a�E��ԝ����m�9���1F*/���f�su��D��A�����T͸�o!�1Yӧ�՗��iN��"?�w�?t8/�vf5���aa}�M0!�ا���9��;��{���a,~$lXM�g@�'���P�f�l��
���#�x��=. bZ����%D�~}�Ԓ6xj��f��ʥ��ʰC�҅~����܂��d|���'f�L��.���8��+��D(˔o���� s�Q��F6��O�N2�$���O��d���h���8X�v�f{�H��!)�
�	���e�Eeo�n_AHe;]�Q�5�v��2ô	8s�1nYm��cK�.�GV_�s������{	ǲ5)U�b���ar�v�9vʄ�n�vܮ�Q�o�p=��e����􋾏*$ړ������}sC�a%�}xI;�n}E۲�;b�.PK�H(N�w��~������[�ꢒ�UjN�0l�v��t�6��	1���}<�iLk���Z��@l}Р"�� %NI㎬cf丫_�Y]5^���`;8�e�
��ٛ�P`�g�<�4C��X���;]�Z��/Z�uBN����O\Q �� �#�$��'�k`��Dfѥ e�JU�����=d9�R43��+���'(щ�܌�yUAG��P���� *Ǣ ƺ`�Meʡ^Y<�#\�&�t�H���Z���Y&��[�^C~G����+�҅ƔC��gڊS ��wah�uF�/{DÎTaq�~ĥ$ �6l���BN-eDZ�w\��C %v
������8j+��7����υ&��N"9WMf�z@��[��yUS���T4�[-E�s�sn��9����`�!���1� s(���N�� ������̏_��6gu��8;���s�7T����ѴH��%� �7�n���Yn���1,x
Η]�� ��`�"�>�h�@J�,'\�/��ҕ����̅2�A-�&�~FL:�Y�����8!�G�5��W�d�'q�i����`^�D�`��qr�[��#)�
�o
Us���-TnQ����tپ�+�@t��~�A)lc�0����m:y����~�"9Z;	e���~�1>�Wz�2���c����W�eE}��-�~��#���]�Y�sfT��߯�LT.15[���hZO��} ��\YO�]��)Q������^���>fr����F���kwƴ���EU��D�%�xRRb��
=?�M���n5�)��,�����|Џ^ɍ�d"�C�1��i�;�(r�Hn53��ͦ�I,�P��(,���3`0�E��
 #u� 8�Fl��":�Ɯim�������:������e� ���m�כ���W;��2�.2�3��S����ܘ!�ܬl��b�f>��$�:^D���N�籗�b���������t��X��`�<_.��F���w~D�8��:�	�]��l���s�����b-t��=���sk�֩
���ÂȤ���yR$�O8?h��&���b��M���H%h���}�����g�C�V`~��YQ�����>�ʿ\�.loU��zK�qd� ���>I3��+���]	�@� P��t�gY32�57O�=���g]�l��*L��嗷�{b��R�7L� /������m�._�L���k���;�]YW�8!_3Z})���I��x��������7N�e+e{�N�ȯ}�`Y���~d���u���/��1�X p��G�Nn���!z_���g\���
;۴����F����IY0X���	��r���l���{��WZ��"U��X�^��fB(��һInO�X�qh_��+��Pc+��;XX�$62`�7`g;�#:8Ǯ{S.اH٦Z=?�&�pj��]r%��a���PI����'S�`�+�LӫA��Q�]��s�ZZ�Q��-�1�~or�(>��ʸ]��Ϭ�RiL�<KJcmF���Ǖs��X����\@GNM����n��J�Q.��mư�%gR,��|���y\P�i�&!D�	�Ԋ��2hDp�T#��
�4�q;`�Z�3�a���Rё����mpF�uF�H�1)Zq���0����>G���n���Z_������
,�B��Wc֞�<K����g�?�i��'CƩ'_��+�-���]�{�x�k�[6��<�<�9^�/?'2,�Y�
�I�aF��$�'��4�ò��8�f�����ar%�����$c|_z�*���g�T�[7��������7�ks,rv�[8SzTǁe�5� c�`�H(��30/�a>�����-k�b��/	k��+��� E�����#T��L4�֪!s���#���9���]BΟۆ`�'+��9ov����[ז
+�9�}:������M�V���C$6��^i��y� ���
�x���]
�Y�W��T������'"4
=}
��n֬�LGd�<1�4�tB1��I&� J&�x+@ZQ�#���qW��Y4���D���W˦�����t*y�����͓�k�C�z���wZ�C�ӾeS1��Ӣ�ʟr�M� ρG&���&��I���)�k��y6����H�|n�T��������U[@	}"3����'U7�3ס�M=o�v�ţ~'"�P�2��(T䯉�E����"�$���K���	�V�H���'��e�[���7(��@Q8Jj��#[,����3YQ��.v�ƞ ���A:h�V9�\}oB5�U��0atWdq���Q�_�3��o��d�Ǎ=�����$e�J��G�>z�x0b��N��ʯ�x��Z��� <��}�l���)�
���R�f�PdԨ3�x��2��r�8b�*�.���P��1vv�l�� A23.�ڜ-��*L{D�����_آw���̱J�H�Q�֡2�t�	�a6�y��勎*p���>��٣�qe��6c�S�BN�5�.kY<p&���_Hy�u��H��֤F	k8�����BC�.���@lh����P�.�yƗ>[w�s�9s;vj�2�㳁�Y��&�~��|�J�b=�[Vg=��H�nk($���M#�u�K��}%@�0{�"ﻃ�;hL8w���tH�9~ź�T�r�3D�,�`"��)C��:d�˪5m=6iW�[�Z��]���k�}=����:pf��-PR��Uy�].��y� #EG�ǥ��^X����uh[6��\�����<�$����h���vP�w��V��u��O$R9�e�҂����9�����v���ʻ��uWB�"{��1ᩮ��1�
�6K�^~�.�F�%Q���(a��v��	Z���Գm6��x���U����(�jش<�}�#��/@�C��w��Q5��������jP�5D��)n6V6g��W
,��?�(����g�6c�q�[UW���0'�K�g���y����|]od]l�d)�c��mݵ:�r�(���FR��q��;���"^N0���d�����h�X�[z6Xyf�vXw���0~��.MW�D�Ub���m�����7�9�>\}j&o42^���I%(����.��#c�2�4NU
�	`�r��ѐ�D,G��[P2=5�����.�y��a:
e�����qA�X���8�*GԔr 끩Z[1�o.=�,���Gj�7,����͙��ZcQ_!.�&��$��>��%=�A+tŚH���Ks͵�z���C����H�@�Nݗ����*:z,�t逿����y=����Ng����XQ��m��m��!��U�����8�c�dy��?xg��\�x.�|?^d��B�m5-�5o�J�����A�`1>"�������������e��oX�lkx�Ż�q���Fa���?�ԛK�T���o�!��W��Z�4 rʟ��lN+	��n�aý�zc9����74{�����}���D�i\u%����חۛk/�~����7�=����s��Pb�xP��V���,_}ur&�t��9�|_�F��Q�oJ8![��S��̯%����tqkG}S\\����Ģ�9�7��<�`!���{��u�Ib�O���=;S�8Ē�Oj4Ҹ�������+�Z���u'�L�а���u�c7�\����uşڮ�<D��&��!�`�b����&�n$���fS{q��h?�x��A_�3Z��4)���K�w���	Fz�����{r��R�j,K����C�`X�Ҏ2��i�ފ����l.w7�����8�-��YP,q8@ǯ�O� 
��=��Z�{���9O��!5h�������@�|���"<޺Kk��i��i��?0�zS�o�O/y��X)/�� �g�j�ߎZ<;�l�u�TL/�o#��Ms�Q��v+`|�a�&���{1�����L��������Νc�����A�0��g�&�Cu-$�C��0˷&Ƃ۩���l^���,�|����qYr��XSC 0������/��;�^i�U�6���%���A��BV����Y싱�gH����YbԵ~z�����\q�����}�1��z���6U����ۡ
�xHbI��r�]����[�6Q<��L�����ܫ����R�v"
l�^��45�/ʱ����d.�`P�X�=~��Y�^���v��8�����l`���(�
̇o(� !~#)���5��'y�����L�z���O�v{q� :#��65wcޭd�&�����Ɠ�pm '�7������TtZU P�h��`���Z½}\4y�Y�������%C���E���8R,�Yz�b�H���Qc�c�z(?����?5]��nR��r����a�����<�#�x6A+q\���i��#R�4i�z0D'��w���\�dA�D G�f�*�(��&��"}��h� ��{bo���'����(\��y n�� �O: ���"�Hu�}�M�檩?1m��]ݷu�y9	Y�K�s�p�oQv:�qH�m�B�em��w�?�p�(�(����c,��e�\����,���	��F�"��f��6B�����al/F}�c�	`8L�<tf�r�~�H�`{���S�Wbb�������4��?+iG����wD{Hz3�أ([L{�RtX"�=�e��-_�`�̓,���(C�HRf��Ye<��o����؈�ʒ��Ч~@Σ�`����#1�GZ��+X�UJ�J���Q}�J��&@�֢������Q�12�М����eؤv��J����r�I�^&���
jx*���:���*j]�jv�b$c�S��̡�zzc!U��=Hݤ3��»��3Ny��������mkf4�mf,?��m�
)�mX���OX�.�UE�

,�I[s뽐F�Yl�&a�������"+>pbl'��1]�p)�����pؤX�D@����^�/�������϶T���`��UM@Q�g("8��,��h"P��6��J��	ow+���*��;���S�UA�2��Bs�c7n<��ۮ��k�:݊ky��=`��)X:�^w�5�����=�����<M�er����3��3s>����}�X�^�M�y��Y��	���sQ��	��@qT�?�q:)tY��W�Y�>U߱C�K:{��w��ү�D���^1�*<��:S��_��Tm���'b�=�,��n��Ĵa�V�_�Ȥat;o�(kY�����Z�o�*:��M��@������&x�Bd�566i)b1���=�	F�Ȕ�y�R$�_3��6ZOHGr�2��E�0S3v$�:p�/���R�Q��T��Uݍ�r��6���ސ0?ar��E���5��ZR��N��n����[	��/�,�V���x�\�C�Y�k¿��1�&q�NVvąB�k�Ӷ����w��c-��%! �O����c�����m������2>K%�X��o��m[�j���`K+QZŃǕ�YCgFK�:�I|�F�%oY�/��g���z���T���7�w�?i�ƿ�UX��|?H��g�s%�6��&WY�����Sjn<\��"L��j���ѣ�EZGYQl�R:to��k����CN�2�rvQ�"�%ni��cm)���⑬U�GS�0�ݣD�67+��g]F�gV���͎ ȣ�}D4�5T��yBЙM���6F���H�H���pcw9u�U��Bn{�T�Cڶ������>8���_YHߎt'�G��łI�m����i5��"��vfXV:�BJ�NzuXӒ��q��GL��l���'���wӹ)��r�G4�����/-[�e
i����&�����~�PC��VD��_c����z���	�|l8.�'��B�2�[;	(��	τ�(a8h��h��fi	
�KX�e�\J_��[�l�-拌��.@f���G�+a<��O9�qT�0|��V�A��e�/o%��S!���<hò�;�F䲈���Z�P��E����T��3}�b���u��?�\L�8�&O���]�������II��<��akk�u�"J�0���P��`�-_��v�M.#�����NK5�#H������X�j%��ω3�#4��z3�~T:>uZ�((P�.���=�Q�������]�����w�����OŦ���@���)�W_&'����Af�;��G+�ձ��Yw}�W�p-�q#ײ��0X��V>9p0S*v�J�$�e��}�&0�9��k.���L�jص=6�o`��p���7�|���2A�}�3�!�3l~��[�G�,���'E�Idv�-UH��Ws�ëe�3�����	��g�0���`b�y����B�U�����EY�V�wQm���s���+P��(_������ςy�21���9��'��4���������-��8f�n4j7d Yz�*��7{J����`'i+;~�YkiS���:�D;�O��\����'�L#CE��?k�q[x b�3l�0��QBlU���yćHt�H\���4s���ce��~b��4�$��ժ���V����).�Ul�n+���-z.�Mf��Ԉ�#�����<��e����C'1=�����:�<x��lv��)\nV���1��\�Jk��8 e�M#�dݮ���I>��M�e̋^=궁�v����H��կ�~e�݊�Ƭů��!��.�l<�#S�QM��u��vg�=ό��;V1RA SL#s�\g�CC���`_L�j�Z�|_oj�21F����(����o�v6�����e�@��7x%w	(!�r�����^�c�%��r.�P����2b$ �q�2�s�3��Յl%�H���\<����~U��� ����˪��{�iM��γ�Ro\)k��N��<�L�%j?�<���(զ�Y;��M;W�f�Ku4���q����>���,�M�E�l~P�x" ���v�f[6`�i!�78�P��ş�4')ԧ��̇ߘc��>�mH���nf��\j� ���?����\���ҙ	�0C�m�ޮ��0&X���*�81���͍��*xP`I[�9#,��>.u�9�'$f"�A���u��Y|	���X t�qnO�_��s�Wp&�d��ɚ��*d
3)��_4҇Ճ1�u��G�X��h��.��$�M�q�L��&�>� �
�zm�D'�2�3�<YB�!w��\E��7R�8r�$�0�y{c�J�'JW���qlq���[e�O=�@��te��kC*��T0�k��@^�R~�w������H��ҵ�0_�Na�^%?��O�L��n�5��2f�Ȁ��Gt�D���"�02]w$�+�A��J�u-?�Zhz�����0t���y��Q4y�~vT�`oQL)��ymS�Ғج��]#EwvO��#�H���<�H�߭�C�1�@���W�ܫ�:�ߡR�:���F
���E$9F��p�9!��Lgg������v_���>��Q�_���%�m\��R�Gy�23Ϫ���(~`��� F �:��G	د����ͪ�~C��e�Ҩ��O�"Ʒ���cƪ%���nf�J�'�7��/:�/����s,��,iӟ~S¶�LS�d�����W�`��U�9I)M�d$n�0��>�;t�`�+8Yr��~�ub��ov��"�L��Xh�g�<��Ŭ�@���l�>�e�uq&����6|B������؎Eh�a���zH�+v�9�W�'��v<-/�����+�����mk�d�%��N;��=D��A6�%0�巧eLUq��r,P��ua)��?\�|E�����$7�3��5��x��@�C/?��굌�V���%���RI�.<�Ҿ���@�������A
���r{˕RN'�V/��� t͙�?-�]��ߞ�CΌ�0��҈Ɲ�/U��͐|7�a�z�\��Z蚊J:vc"r��JPa���G��b:�M�+P��lv����\yU��-��E���|�����-p�p;��8�B�Y"�Vsy�R>3� ������k<}"�/aDsp��N����F+q���T���.� W�7	���FE���ľv	��$]�ٔ�f�Θ\6�mh#�ܽ�q��f��Z���hѨy&�l��613�}���F�L��(Ms3uX��ڲUB�$�Q0�@��F, /��:����)�G�8XaH9cUe���}C�����&��O�bz�������|�E��_GC*������u-c
=��\�9˃6�����ू6�>�z�
e��XJ��T�MM��,؇e[���*��1���/�8���7��P'}Z3���c�D������'ϱ�����$q[D s�s�N�U��{��ڵ���֪����%P�U�2N'��o[�f���I��q�و?������h:����j��3P�E�t����g�8����E���	�+k~�G��4V���>�
�W��%�k=e�y�v���p(1�?��P4��:?w8�q1v�+kjo�R'y�a~���&�+�� �J�mG��ϡXḜL� l�v�M�M�K�"NC�����-�<ʖH�5o�H�v�i�t����UIz!%�ADp]J�\��W��Op�,.�Dl�?���,�s�,��g$�x�||��6z��OX��B^u���#��>�q c�ͼ
dg��P�Q����F���'<9�,>�C,�8y�0Z���XiP���),�iJ�Ξ[�X�Ɨ�՛��Ќk�#����
���[LD7���l>�ɳ�$��3����U9Yݿ~�S���+C����d�B���UU�G��l��� �F���KJl������,z&�;�._J�G����I����d5���D:}�+��d!)A���$�񥎆��*h��E�
>rq�݂Friu�&eI��;�n~7#�xRs���p�u'�h�Pob2 ��q��u��=Iȶ�p�>ڑ�?�k�)��`������R�g��C/�]!,T�-_��N���_�l�y��������Z�����l���h����YLU�����(ɻ�ϥ��[��
��MkA=;�[���}?���&t��U|��R�����6�t��. �/�j�;@	���a� ��o-f��#����)�� s�O�wt�t�KU>[�m�{O�D��w/���
��Ry�O���Z؈����!�"�O���Ko%������cۘ4-@�Z*�JoZ��-����)�wP�;�wy\lZ�^I��ǌ���71dZ��3�J�5��{O�W�2�gqT��~i.>����8Ķ3w��������Tn��F~�X%50h	�4�i0���h�	�����5=I��=�#A��T%y�e�ä��U�myb<�u�;�����'���faQj�m�	Oϋ�b
^��8�Xct�T���W��UdS0e�yVh"^�_3����&W�G�u}W���ER���s� ��G��,��uN�V�[D
�Y��!�Ǉ��F�T~�PKq8����C'� �Q3�����*�dRl�<�`D�aS�Q Y'������0ծ��w�П�sNi��d�O�sF�-�^�z��I����R��8`�nj����ԗ��.m��W�58�0�i�E{��|������Q��JO<�j���ℾ���6�P�V�a]ҷ����8v`��A;��F`}�]���L�^�^�Z@L�k��y�a��u�Mv����h;����m������.]ѣ#r��a%����M_�R���Lɉ�J��[*��r�'��ȇ�H�!>/Y6�޻�)��q��EY?�Ɔ��*��%'ȡ*�CN ��3f��/E!L5��C^�Sy>�hբ�U�Vi��,_������1�q�|C��[�E�d�pY����5�k�L�9�Y� �3����h� iˉ0���׌%���U@6��38EJ���(��/˪`���M��w7�����*!����6����h]}0�� W���������{��(�PV�U:ɹQ�y
��Ot�=$��(������ (&[���镐�Db�9�@��n�;�G�ҺJO��"�E�P*S ��S���1q͆򈙌�?�`���,C%�vO��$�7��5&;r�]wJN�����W��;<ߏ	�Uf^c��F�Q-Խڦ�ףAH����7��y�&��9:gmG�үFɌ�GQ�j:vw e�7a���e�=�^�˜�E�vS�5E�y�wC
d 3��Y	%��E��*�[�%��J���k�!�v9*���;�#f��h6J�ة|�)�.&�Y�,��O
������Hv#3Sk%I�ec���^Z�枒:�E��~h���j�2��=���on�#��l�t5<�K(�S��h�l%����'<�U�:Tx>I[LP�qP����F(9�{��Q)���;lph�`�G
�Q0�TUN�NBs�)#�L��|ő�#ʤYc�.���δR
��	inB����hw1o�
��{�أ���W�Í~5p`H�}�0�̵*�ntYr���^*�Q8m�)\��s)uMp|�������g���bBb�2yn^��5ts�P�5���y_m6g��Z����d�>��l#�w��ׇH�ѹ����]׫h�y�:k}��=;��.r�����.���sZr�32N�\cbw1����\h��.�ov)����3��D���'����,�^�<G�%����d�L���A�w?p��6��v�oSҦ�	*V�)�0V�\-l/���������t�/7�\zSc�2S�#��������7]\��S���z"{�N~�-l��"�;%��Q`�cM�8��`s���"�/ �QYi�s%Z�T��ʩ�.~�A�(ᓥ��ne�j��p��{B��>�������/gM%����
����#.����Y0g�{D�V_u�5��]�8��͚���p�x�z7G�5�ԅ�����m'.p���9�x��`%�=N����bV��2Ų�1�=NS�oG� �����N�ت�XН�s�O�����=�119��|�5���I�OЗ��9�._����2�֗	8�\������E���u60���0��X��U���9/芥DU���*gY2�B���=Y�Ę4V>�\�x��>�����D/=ŀ����lks�U��5��}���-v���R�~A�fb��W�1O�I�2���J�F�N!+��8�?���˹0:�V7]�Qb�ƣ{���Em8K��^B�h������oӖڈJ��,Æ8���P�=m���f�W�zcK8i,
�n����J��~��G X��m��Ko���k }��n���9Z>�L�Shw��+xV�r,(�4`�B��?,y޺O�*���N�/�BV���}v��o������M���6����բ,����Y�b��O�>��T<��75��G�c�k��~��Y0���8��s�up��ir�+њ+��ؚ��mY�9�v�8��0�=Oߊ7ʞ�>���2���r��%��y~G5�X��1�6�����&}�|�`=e���w�P����j�t;�a���^0��S ����0RE5ʇ͕�4���u'�+kM��|��eV�&ݶURDJgᐑ�Ez��>>��ߊ����qs)�� ��, �����[ڣ� T0[~����Ki�_ȓ߬/ܦ|�1�:_� ] D�JRK�������O���������w��:4;l��sp�]�Z[��)aM�ܧ�5�|3P��<�-��h6���0���Oޟ$���)������<���߱hv�q�ɐ]��Q.NM[fHQ�'�IwH=E6�hȘ�A�ҙ^%Tu�v-jWp�����I�%kk����'�d�K�+W��vub9�3 6)+�3;<��ǯ�E@�/>���gek0�&"��׋�<wY,���"U�j��R�[ޛ��S�q�wn��x��hS�'
t�!+�={x�萎�h��g&1'��҄�jG)��As�b@��.��u��v�U �wV_�B`��~��(oN�I�׆f�	��U���U�w��P��U��孢d;����X����+���k�G�%�������?-��#cYD�̏����d�q��g�4��L:��Z��o��
r�jf���AAd�+UP^$��*+i���M���y�f��:��r�����sH�f��f{��Q��Yę��D7����.��қ��"p�Ph��)ԥt�tEIA��ĉ�:R˧0�&6ۢuO�a$1˶�$ԗ�	P�%"*�L��ܶ���h'1�����n�3����Kv��w(,�����B���Y)�I����8���>��w�/�$�-9kc�Chd)3k���,5?��[�E������]`A�1�֭2笣AtN>�K��
�� +7�F�D��p�,.(1�z� u ��������hg#y�I+Oq��������+[��J@�����jl��	����iV�.���� \�W=�Gn��(ix���eա��Wu��)�f48�?��ӯ\�.��t�(�0��{��󥔯���o�u���˸� ��7M/R�h������+�Q�G pw~�ow�c����k�rl�>Pk,���K�ѯw��(��~������g��YJz�|'@��ۈ+.b���^g��zD�a�p�z0�>�[��8���t�jg k�A�Z�g}���eI6�{ր�b54���Z�b��I&qZ���1�I�}j�����Zl6�g�"$���C���m�D=^�����M�_�)�o��X\oJ����w�B��{���)5�0nކD����a<=E����i��	�dl�Y�N�����,��&!*�UB_x�d{1��旇�Z�*���{����C?�����w9�bvr���;c�q�	��ֲ�M����q䐻\0M�QG�%�;�K��.^���*z&�;�>~����&@܍�%ظD3{��?��/�S:��E�ߙS/��G�A��<��ĄtA:�_5V�Q�K#�2f�d ǂ������]�?�|z7)Lo��5~��Cz��M��g��F �� �#.l=S8<��5W���z�MŴ�^�Q l������4J��*�H>�2��w��n�k~�>�$a"f~�S5����ϟ��3���a�3�3��j Dkw��T(G��Hj�8�k�C`&��y�����g�<�w���Ӳ��-z�^`�[p��t��O�����r���_����i�C8��.�W�A�� �#�uA�&i^�t�XY�:�r>�Q�۝7�n��)h��( �И+9	�l ��sd҆̌���t��rf�u^�XDg���N�\��\uء���P�Q;�x���`|g��A��\���fF��v���Uvү*L	�l��j�Zo	7/	C�2�+�H����3@������H�I���6��jh|c37�@(6�~3^�{��\�G�0彿A%���g�Tb���HL�c���~������yK�����N�[���U����LW��6?m�^�-��@`^����Qgy����k|��f{F�o(���߉7�s,y�Fcc�as�^����B���t�Ƥ�]�*Y��N���(�����x��f��n��K8��0���F�y��zN�JkQ��f�0�xmB%ݡyx����x<�n����Pjo �U4��ò�w�RΚ�F;��F��T,\~;W�a�e`�h^��L0���h�B�A@$x�7�� �].1���6�3ϟ���5���/�����FY�
��W��'�0�}U����Z<�L�݊o�`�����'d�9���=�R�#�� ��].g߱d*n�6���;l��c�2����J������%��]K�X���h��}���z�]A^�jQ�5����0�9��U���B����W��1��W>(��.(<`���BX��#�}�h���%�-u����#b��wX�Mzz�f/��"8�Y���&(d^j��+_�Y�
���(�a�{� �D�ŧ��H�aT�P�S#<�(�b�<���1���-�?�����V�z|-�����w�M�sƓS]A��} �s.k"�o�l��{�����ܨ�V��9�8�x�ށ�3�w� �m:�Jx� �m��F�g/,ܞ1wM�Z�g ��`c�$���t.aX������|����S��\�l�Xuz����q:rw�u�v���λ�1��w�.0p>�/R���E�	G�sOA�g���a2�0n���ӎ���^����Ry�y���
!���	f�x`
�}��X�j%At�M�]��B2f��*�תj���4�t��}�
��\��i�(�cUz�1�%ΟU6g����[j���j��>sHE���.9�-)}y �~e���ʞ��\V�~�b��d=��@\}��y�#�_��շaE5X{iÍ��K9q�qC\-���S�	�a��lRX'��c��Q����@t������-��{&�V�%���Zo��*2ext����)�nn���YZ����^��:~̋$&�C>�}���(\��P�8�z�+�+�&�k��� ��T�~�L@���k���%�:A����$h���`1>/��X�Q��m�G� N���D��"�߃�9Oa`4�=A������#��r��7���[Z���]h��3!�j��
�Ϟe�vG�\<i�3��5\�ߊL�h@i��i��b��ֲ��m?Ouٌ#���>�K+����®N`<��;_���ѾX��y@���M�T0�I&�?B�7�c���i���!��H	�<��.hM��G+-�}c(����ʢ�`f�������|~@9_����#������{���B0{hq�[KN�b>���Ĩ-
3��vRs�Nz�I}�*:�f(�m����,Z�ֆ;�a*
�n�� �]C�F$�"�*�_�C���">z�jv��6vX������5�]ۥ%�� N�Q����$vt�gz!N|�"��5N&�7���yQ0.��$L{�P�ho1�7����V%�@p:�jM��^�_��Mp1FW���"�����r3d�8��`�E*��@Q,_�h���o�n%,���\DH�E�Վ�a�NV5���-���7�@YQn�C�?A��X�V��e�A^q�O/�Ѫ�P���V?zXp���O�:ɿ$q�,JlH�Z�2hg��>��4���-����N}�%W��E�����h�A��o�ۍ7�2�,�ɶ�H�.�Vmk%�zɡX"�N����0絾�]E2���%����Ud�Q	����8E�ب�ӷ#VOE�)s������Ƴ���~
�0@�󭬗� .V��H+��	���phƒ`��
k�ɏ�F%q�'&��JO�w�}�\������4�-=o��4�D�!���nz����깍v~���P�k��pj�;���J�d�޼����?��֮�*[]MTϵ�T�%������D9���֯�����5nM�!0����9��9��W���q�)���s4������B9X�i|��5A�9��4�?+��;��[T/��ܷ�ť�\h�B��D*���+8��Q0���� �%nN�Zc_�LL�X,k��eU��lƲs M����(�RԻ|ۦ��+��+!���37�?5�
,Ҹh�r�vR�i��43��xm������F���}Z	�L)긺�	r������Cd0�(u��o[�������:�U��ˬ�C�X���'=�C�'���g�*�(� =S~'������)�h*.�-��N;��Ǎ|�<�k"�,,d��Z&_�O����/�Ź"E��X�e����������ZBǵ�[K̜��_�=�#��Ti��C*���˓~�5���,F�"ه
_V�1<M�YP��R��-�f�ȣm�Ќ��s�oe�mLe���;�k([�&� _W���ɘf���Ʒ  <@�}z�x瓚�	�ݿ�H�rG ������q�iUD(�4,<X��}��~�ݹ�(��Nƻc^�����C��� Xh~�ׁٙыp*���� g\X�$��q�.���-B~6�#����sO$W!=D�}�(^[��$�&m����>�!}���f��%Pq�\�cP��p6o3�<�4cޤ~���l�K���o����լ��hf�����t["����)k;�����j��`�XY|�!��������JQ?>�0%��@���������$~��R[)	h���m!8#+��nB�z&���[��u��Tph;�/E������-����z��K"a3���%p׺���MY"nLN�_�<,J��b+�s�o��n��' a�1�	ᦞ�'�����ދ�m	
�Vx�UIs#:�I�i��XR0��G��0�jaR=��w  �wD�4�:�K�N=��n��8��N�f�#��]��������a�Hq�i�2Pv��$9&\j`�A֞{:k�%[LŢ9u;���ߕH\ha��H|�6���{�&A�EC�c��{T�UI���v�� ��Q�*�;@�J�:./�)������pA�?�F���n��jˆ:�P��i�f��eTҌR��!;sn�}օC�Ҝ�nG<=[wl�����Hi�@g<�"S/�?rL);��G���g����ُZBK3�T��f��a`�)t���Bh�i�7)７̫&AN]���� ����T��$�CD� �-ط*u�~��o�?��^m��Qz��oF �Q�+�e��ƌ�.��Z!7�8d�J?wz!:���M�`��?Mf
$��x���Hں���~�IMe���ƪV/��&[�}�yy�c���p����h�F�1q�>�<,=5�j/+�4G�Ti�H��k��*��:k�� ��t���5���`�큧�U}�c����C�G8���k�^a"�-�:;r�tI�&��1]]�ۇ���4Tͷ���Ǐ�T��я'�a"�A��NG#n�0���T�BoWY��ۄ��{UZ��*�s��e0G��;![|��ݕZ��2��������]O��r�1G{��F�TZ5����7�ˀٕ_���L��q��P�WQ�V3o|��i���Ii[<�h��8��H�~ RK�)YQ�8CNߺ����ؔ~��5�d�y*��u�|x�B���\`(V�������A��ulT�����f����հ����i���DkFt�����|g�4<�9�N[���� o��r���Q�Q� �%}��.�Lwj�VElGY����H�V�茖}��1��,���9����:����R�Os�kn��V�7<E!�q9�e|ֳ�sV���2q���䒺�v�vj>H�+�8�
<��Yz�Gm�pYhET��b ��h��"u X�U��E�[�}�*(\��'�Jp~��D���ƺ�R4��<s
��Kh5���y�c������8H���J�F�ZĨY=Y.2y�2�)�'�]�^gIR�a�M!$���!t��#�H6O��S��V����F=��ϑ����C0WT�̼@fC��>�ML9O��aji�Q�N��-�.����J		ˆV��g4�Z6�z�_^����Z�Y�4\`Ԅh�&ET�sBO����I��:�E@s����ꏩ����U(�n���cS�֠nV���Od��M�_#�+#�t��7ԍ{�^�n��h�P��(i�W��AD�K�f~�0�ヱե5ߋFڃY��&r]q?�J��Y�db��2��`+m>�Wd���gzK���A�k��˿�g��C���~�˿eL�h�|y�] �m���}>8FR��썮c��/�H[
-������j�aH	��~���pW��l�̉��J�e�P��}��+9`ǡ
(sj�^�/# �:Ib�rm9�׹2��b$�R��)?.�>p�Q��1dCcyܙ���6�Ɲ�E0-�]G� ��qEץ\v�w��S��Ӭ�s�
3��
Ѱf6�#�q�U� �����U
{K��!�^ko���du���7�����K��.�b�B�?5uT��4��n+�+&z�_/�NХ.\�dR������P�N H�����k>���X�l��C�Ҫ1e������A��^�t �R�t��܎n/ye��n���#\����o�+���iy��E��uu4�N.[����Z;'5����	�֡Z��`!.�}��&�"��e5��I� :A�|ߒY��V��VSkޫ���X7��[MA��E��ј6S�چz�܊��K�5�'L���]̈́&4��I��4�s� `�Q�eb�*!C=�'J��}�?1̦[Q}|k�6�:�m�+�C�"�0�;p9�h�B&��b|��?	���gX�^��#�����N��Mu8h�t�p�Ӽ��e�	r�G�T|T��!�q{��ۭE|a����(�bPF�� �o(��ĳ�2c|9���,�Όfb忖���BtF����M��?�.&q�-/�	��7��ԁ�Fj;.6jq}A��"qO�dT �H��܊�p�Z�=�
Χ)X �¦��(r�Dq�4U}���-��v�X�2{j3��د^�$���/u'�d~^�.�-�:����(g�q0���u'"����-�,D9��I�vd�;��^H^Z|�������L��٩gpN�[k��O��d:}������BzJf@�d_Ty�Nq�w���H��)�a!���I(o^�O;����u��Ś, ��Vv*�˨X*G�"�Z����=v�����v�������4��/�4"����
LTYY�M{�L��X���yF��4�/��`
���
:�wݷ[���~��F�9�wU��Ӄ�����������F:��>l=B?l)c�^��� ���"b��8��8���)����*S�e7^�����Ƌ�x��i舦�6��3L�쀹_�~��P�����E���$�^?6eu�nA���n�5��a��s�5����~H�L�@�oں NS��y�?�f���d'��H����X#�����o�Z�3�ϔyF
����@�zs��9|� �"F���m�sI�5ٷ˚���"���N"�o#[N�P��7Ǵ���S��l�I��n|�R�� �AbTz��e�1����5�W��_�\"M~�<`-Pʲ�U]����A��;���`hQ�R�����Ǿ]��M�����4[dQPU;��[J9�*e�j*�E�y��5��ǡ- s�?Ռ�R��;�v�l�dH�2�g5�4��]BHכ��������"�uy�6[H3����U�ʳX�V�#�	�I L������UW���4 �m��+�xݲ�@��&�,b��$�Rp���E�)�q2��l���1�<M�x��o�&b�v����s�=�2] ���.n~s�#z�#��ѥꖛ{r��� \q��� {��Y�G �o������R�5�8�C:s]��!"ǳ��V��ĭ�8dRn�bԸ��~�	��D��,�~MKI�+5&x�%YYj�L�,�0e7~� �V���s���?�g&:��8_P0�5;)t#_�]}2���E��r�֐*1!&b�a7�I�C�sP��h�)2L+��q��b����$�Q��s�X\C�e$�
����R��(�ȟ�H5?���){њ�F�#�*q��~C�}>�B�^�i�Ù$�[ 2m��A'���d�"5]x�:k��Ƒ�@^z]r������B��Va٫�h��&D��cwɸ���u�ਗ਼Y���Ʀ��D���I��	�o�hn�O�(L����$M��oD0t綆� ��?�? F[dak��wKaK>�z�J�Zi9���B4��E�Z��O;�n2T f?��*�|��q�H��g�)zu�|�L�x�d�
7�Z�,7���)���װ���P����
�!��%S4�4��9��0{S����1�Kײ��=���J���_2dUS�I��{bx��޺7����P�1k��ȉbX�O��Ϲ��� �M~ϓ�һ`|�¦Z��W;���U74㑇���T��3wi�H�,��jl��WZ�|ꪳ��)[᝺���&��I��N�	�,KIU����A�^�/v@�d�,��k��粲��B[��-I�b%���}Q2�N��?ҮDo��ؓ�Z�=�����y�����o(�B�%�nEz��	�aH���[�"(N��d��NW�*"��O�O�� }}�l�F�;Ɓ��>���H3�{���a��@��~�GJ�;]A����k����1�= �%vŌ�4�y.�Re/j�l�M�~�z9 &����/�PD���6I�O��i?x�@���<Xu��:�U.��&�;]E�;�q��-T�2�`�a-�����F��=���H%̋i0Ih1�Ԅ���i�\��I�'	�������Q���.�z����/�w�B1�c�|(w8V=�]�M��^{D���?�!��Htc�0���G�>�繳5�K۫��p�5��$�k�%�����5���N��$�ؿڼC�-���2Ud]�^������b��53wO�!�mTW��!鱋R��ԯ�g���q��F8Ҧ�&-_j��&�/,����N�n��|���G�����׻0�N�$Ɇ�]R�׈� �
�"�)O���Bm�&�`lR��tc&:�>����7�_ͯ-�?'�s�P�Ru�<�G��S�(.�k2>�9�I�$ܱ�P9�p�<��a�1#���뤸xGry�0qɿ�w�65>�,��X��O��R n�:��Qf�� /C����F�O ?}jY� j=�q<���و%v��T$�M�PK�5 $8�ӡ�\��TG�A��_����aOC	��áa��(ѡ��v��*۰�m�t"���GEϓ/�1a���=�a��]�K���F�3�k��x-o�e��-� ��l7���
]9r;��.�e�����$�ڞV�yl=G�c4~��5T�!�B���ѽ�x:��c֏�v-�"�p(j��e�*��4��/�B��~7����Ͳ^���u{��]�&+�,�QY[��>��1�m!=�p^��#�	K���$7|�˹�#�����u��@��o3���/lM��;}Q�ǎ;`���G�1�vak�c�L��������$ю�^�}�φz�bZ��W�p��uLK�T�6K���m�1�'Nf,r���\��>)�h(���� �y)�3�1&ʛ�";�뵷i��`����j�������U��� ��)�p��T��Gr�z����% �p:5���[�QK�q/�zu�ו}G)J�5<��L9��΂=
Q���Fg�~9�N�"F�Xk��Ϋg߰��CG;m��0%�����n�Ȗ�,�0���e�|���ٴ�/1m�:|V�ޯ���>���7��� �"δ�N���#�ɳt~���2�����sn�����KL��n�2d��)�Ñ$6�jS;G/��1x�OH�TC߉c-�b�~��W%��	Z��e�CE��8����"D�`����L�P	n�[�?�ß��z���0Y������x��\�,�6q��+i���Dd�#�PY�h�?V̂�ڠ���,36�x�5���ؑ��1ExOdk�L�}�wͫ�W^����)z�38Ξ�����\*�K"��{��?Z3�!pε|iF�	�.'�c��Z=C��� Q����1��8"1��s�q ��"W"���%�Ҍ�߱�5:��j#N+q�.�v/m\ި���v3�%�u����os�<���:?��bF���-k���v�xXt���e;h��:|���-�>�@����u�E R*�̞|����{�	�_{��cE0��� k��Z����z�7���u�}�� ������cM,�F�f���:��s҃l��|�>���zrh��ܣ���͚:��ǁ�F��Ӧ|��/����j&7N:���`�?�Ux�����=�}�6�%�pt��ր�w�.��h+ςlSA�ZM�穗�a�m�9T�^qB�>P8�͊y�Ԏg,��SG��Q��+��]&� �~���`%=��^D��_,��c;���j�P�����;z$�M�����N5dvRI�_(�X�Cr~�m����ͤ��g��S�4|3!V�3��s�*�o�s���x����|W����*��S�B@��C� �#Y��d-���s�모_��!]xy����$���ΆmȮ�-w�@1�X�@ʣ�:�4��/tRk���Q���W�Yh����ŸM����`f�F�Һ^$�n����x���:�	P�0�$�s�� ϯ���y�A�\(q"U�)-�/�*�;`v4OE֬�Qr��x� ͂�r��6�i�%.';���b
�Y�� �o�(4���_����:����E7�Ld�u�寐����d#��4����5�N�m�j�7���( ���v9i�	ɾ��m}��v��n�[T�H�n����?b��4�Œ���,��-��6���!����D��vC����P��ȿ�?�8Ai���&p��O\�P�fݓ1Ó�^��7yR�i��V�tb���=��D�!>ngъ)e2,�}8r�᫥���
��b��Oc�2��oϠ#��Y�m3o�{o��1`ų�-NU�L�<Y����l/$x�#�q(t��&�݆��Y�����| �j܈�U��q���G��U���3�1��V-T��������/�_3u�؟+KfB�#8_[��{�W6΢1�'��(@R��YM�&�������H��-���kZ.��I��pBF�"�<_h�G���O��z��<cr�����#��1�� t�=	��m�3��e��'Bz���h�ׯkο�Md�8�� �� �M�+�=٩1���S��% �Y�0H�TJ�Qǧ#��mv�*���_7h� �Mƻ����7�-, -���J�&��"�T;�mݳO�����d;��=���!���Yt�F�7g̪zϥj>��X�-m1�#~�*t)\�5>�r��H�\ͨ��@|k&��k����/����?O�m^�?��we߭ц�	�.A�uL:���}�ͩh�T�tY�Z�������V�}�Q���r�C:�O*��ː4Jʮ����c\����â�8�J��st�_��Y��T��1��xr:%�Wne�؋e�t�{]�p�~;���<li�sJg�P��R�!aY؍`;o�ڥ �_��w�p�"ڊ;iX��LKɴ���R�<v�4�n6š�� ��<�`��S��xi5����b\�?㭺G�z�%�5Z8���d�m��U�E$���������,��_ѣ`@N�sxaK����mb݃�+��[���)���L
�c�&:jO�J��5��JoB�,d��G{+P����8�2Xſ��n����@�ڍ���:�稼�s�m��->R���H,*VIe9�=�9"�Ow�����E�5v�[���3(�@ck�KgM�L�L�����a-6�\/���^�U��p�y���i��Ŵ�Ǆ1��H|���tL�%�h"��E���|-���xx�#���~���m�ހm���yt��?�l�ޒN8�ѴAd�RǽʴϹT|�-Q*5&fl���1�y�"���T��.��� ���5h���O0'����$		;nz�L����������]g����L��Sa��fGy�z�������U����n@S�y�?u��"n��I��~2�@U�։N�g+�Bmߓ����(�{8�$�>��xF��(����1Q��
;u���*|T���ԩ>��Sau��ю��.��r�xxf%��Fm{_��9!�n��r
z�2;�4�U�nE���[Vu����U�,)�i��,�ٓ�%D�T�E�t�*�e����%7�f���Z��[}|�!�A�:)���v�`�p���{}��")+��v%�nX�J��K���%tjK\�	_e�ϳ��o"�bxvʖK����qS?���|Ҿ|�S\� Zҫ����j����қ���w6J���g�?����Z�b�\@H;+�{Nq.���(TQ[89�q�רC�Ղ�k#��t!)�IܪG�su�\(��<������q,�����4���2��1��l��we���W��f��Z��F	۠0�������¯I�n����������0��:Û1eό$�\	���7�xO�!N�f���~vf�j=���Ѳ���(w��)1���É�x�!�G��W�R);*`>%�I����%'VbYy	�EZ.e���x]s'� Ȥ]� �ҥ;��f��vb���7~{]�z/Ai;�:����XZ�`�y������[3-�z[�zp[l�9~1(a���ڛb,�g��x��o�	6�w����{��b~Q�o@��(�5' }%���Bg���c�cc���~tq����&O�������:^��<�bϮ�.<A2����()d%��6���t-gEU ��%��՘7�r��O�fl��1 ަ:���S�k2}��R�<M��_�O�b�]��N��NdW#�T�޿�qpXwus�ч9n�C���<ZMG�B�ɺ��В2�ј��@�����l2�~��t���P��\�IxlF����z���iU��~8�\�������*r�U
�A�v�Ң�5��K��HD�6�Ǐʇ ���w�Qu�cU!}�\˲���V�r����V�0��I2�E�h->����p��e�� ��V��o��nc��q@��bed9��\Ya���-�jJ�s=�(���4�JF+Xʗj�H�/�d�&������Yùs���eMa
^�n�Ӆ��n���ITM������W�4�u�tX��D�	}�q����N�'&hwp�kY�W�a�r�ڐUk����*���a|�4�9�(�N�H�C]�ى�;���+� B%�]BB��>`L�c�+E��� ��(E�%Yï�FW������� W'���5=�9x|���c
�
�mTwz[<�����GP4�����_rQj	}8xQ���>*�%9�##F��lt�#ε�@>x$tn0���I�W���$`���.��}�gyԃW��9��Sr�A֚�\+{1�#+V�ңt�"���(�\؍�g5��(U���uDW�ގpK���2i��%���6��;y=�"K�C�=3Ox���E� �: sY��KTǑ��ʡE���r�Ϊ� ��ҕt�<xA���qS�04��'� �h�$Tc<��tn�] O���I�?H�s�[��2È��~�xA�}ŮM��V��S����ѮO$]�썘�>�,Ԫzɽ`K�]蛳u���� ��Ӫ�z�g^�Ĺ���޽�����<�	�cw���&O#��
p!�S��z��;y
���h)�]v���K����VP}�X��؆^�xa�j��Z4�=6�+W*ZJ��k�.��W�4�Ȱ�B��7�Lpy��Ws��;N�m%e,T��I֕q-{�1��aU�l�w����%-���f,7j-�C�&�Io��$c7���HZ6�0��r`�����/��9��xg�Fm�T�9�v?�;�4��3?{�%��BVI�t�%D�����D���na�2"�fAI�,��@+�����A�㔣ɕ�r�aafُ�2��}����D��wk��3�)�{L�&����@���a��]ŉj�>�R�WA��d�C|wWr�D�)���C�=�"�]��-5
� %>]�@+#
��i��r�<4^y�C��^n{��42M6/�XBy����ET������ y�ߜ�7��Si[ɯD��ݪ�Z��J���z!���t�E�s�N�]���p3?|V�^7+w
��7�n]�NG*3�-_�~�"��	��*��PF�[ ��j��Z��'���q-�+78.��[��BU�;[���#��8��/�5��fK��a2�Z�Z�˟�CjV^Qn^�[^�CxE��U
3�$ᮭ�rB�〽&�B��E�B*�\w5y�������(9i�&"�,R�A�lb�� �J���yCb����l��x$��^��8�c?\���jR/$fN����`��8AOk�6��s�M䘅1�n�ʀaVT�9A(��.�x���K���1W�"��0n��~���&�f�ۍh�#�H���jrr�ht�R3~Ճ=�n�~�f�B[�f�n4�B�O�B���-�ЩqP���S�~1��0"Vݜ�6�!V��6D�r�e�z1>��N�8��0eō�	LG�'��K���#_6��{k({�P�w�e��q��]��J�̮ ��#b�چ돽�&=A�Rbװ��;>)k'����_�e@���;`�?�d���օ�5rzh
	"�Cx�g�Y0�;�M� ��\0����,gub|��Ozx�j=|��l������>1�3[xX5��*�"	����F�Ĳu�»y'����;�y�q ���蜥H�|DtG��ŭ*g�	M���p�Ղ�\6�	����^0�2��2�9�K�t�%�闢y%-2ޘ���c��/�,7yi��A��5�h�Rz�dH�a�'/$za�I�)6SB�lMv�KarM�sc'��P����ٛ(5;$柷0����*�"��{�]��J�KH�1r�u�3[���HO�*	���H����֧u+��FcgO\�&�|T��c�O�OGp�l��y���M=���H�����8A:w�{h�LM�(���
g5e�.B�eaNn� �R�ܛ���0(c�=��l��@{5��l�$MD!?�%��F�b���@��d��&��xTX�R�}\�c�ń��ā�^�c�&]�ő�)p�o _uZ�摳59�_��d���w=�U���i��!N���2���{�XB�d�7&�b����L�GT�y��a>�ʹ_^
ΟV�H2]���.M\�B�l�/]�]�f�LW4�Խŷ�`���'�](XǲTK���"=	����^��Е?�ҤҰP�X;�8�!N�m�69X�/s�̠��G��Uv���c����c�i�[c��֘�fp�Q�1�F�-�e�ú�ߦ���?bt���?f_�l�b�FY^uN�'T���o�i\t�}��l^X���:.kO���BW�l���:�La�0	�h������� �L���\4)&�_���6�y���T��ݢ�:�����Jh���AbDZb��|�����~O��D����!�����Cw��3 	�v+�P���d�8���F�R�E�B�� k������_Eb�y�|)s����ٺ(�MT&�ÎJ�Ql��E�����#,=�3���k0��(�~�ù��rl�E����E!i�����PHr��ض������&��|�Q"gMS��$R� ז�L�c�߿��f�4U��x�Dp8n�z��]��~�u�EoLF]d��c�2��d:����Y���h�Yu[�1 ��挕�؅��B�Էzf�^7�R�'�t��#��ʃ�U�^��� �dL�����؁�Z�0+˲b-B�F7cȕ��h<"��V���5��F�2�L�x\r��nBx_���Q�w�y�����`���kwZ���Vԕ�$�]��m��2c
n���|�|ѳds�Bz�O�2�%d�5�m���N�@IA��B��V�f�(��j��C�+�̳�R=[I�w��꓌w�t�#}��ph�����xY�#�������n�o0���0J+V|2}����*6�LR����C���t�����ߩ���{� �گO{"G���(Y2�hJ]1Q�r?�m�H�rer�K�u�H˅�`#�s��:�^�<Py$�5؜{nھ�|^"H�	ڰr�+�
J��
��*���*�@�Vxj8�W�ZR�� Iwr�������[\l���S�Є�/F�Gm'n�0�[t-ԇ��ڞ�.DODI���=՗�Ѽ;���� S��9��� Q�()��K�J ��P���I)DՄ'�$1�O�'I/�"!�4�c�P��;��G��j>��Ɍ��G�ݩ?���p�;���|O�_%�>B��ne+O�j��[f\����� �E޴���j-�E$gGi�� Ofe�m���g~��N��IY1�����m�9Y�B�Q���|rڷ+��*j+U����5 R�Bz�h����e���"��9ɤ�#�>x��!:y2]*�ma��$Qh�/>"�=�;� ��.�~�ٿ�CgrDWv]>�#z�k҉ý��A{�]� �j��&�<�1�w�f*� ��)0�����	���Q�`.@�7q} ˵Y����[�V��1롴��3�Ol�K�9����
�	���{��8��9r� ������¦�c�CH�1��4�o��U*P��C�R�����#�u�e�������c�-�jΆ�����¶ �W�G���o+ͤ����<���S��2o��h5���y�w\s�1�ݺ�>��Y��Gl�T*N�s�n�sIE�'�ɠyџ������jV)�T
F�GU�� �8��~��o�ov8���AJp���2MidH��J��F\��ȹ�^�cU�$KH+�6�B[��L@Im�D���X�A���r��I����¦�'|�NY��73�b �J_a�L�����{���&=�Ti���_5��uG�_DpW�ϫ'!�A� )BLa���:�8f�>���N,j�P��z}!SE��E()|����=��  ���&oؽsB`����S����5/�2Z"'Tؤ��rl���5ݒN"��}��q����9����j�b��5�������{(,܈��b 뭰%��ʣpF���N��`j:4N�ӆ�v[��MwWd���EH����x.��Pn���r��S�g�7r���+���NI�s�P����;�06-���4�"m����z�;��%E�! ��!��hՠ�x�#�5d�M�ۂf3�Z�v��u$w��B��Ρ��-���{��5>�d����� ^�bN�)d�,�'o�>�W�ىs#���p"��~��� $�D��D��s�ZUb ;�����������?[�<nX��)��r"`���`�Vs=*�8N�Y�����3�p���4~b)#�X���d�4Yk��0��m֬�	qrq�������fg��6����� ��@9=rI�s�?d� �G�`�p|-�gKY��i�&,���܃Am����}6�G{�X7�Z)7�3IWgYb�V�����e���a<IT�f@�v�:�~}���>�l7(� ~#�}��k$QZU1�ʻf���]�E�~+۷���
i%�X���/�m-ba		sU���',��*\��v-�
Xkx���Vѓz%�O����K�q���g9r>)��=�_H���Xwh�)?���F���0��V��Qq^��oEx7Eg�@%�����=�F	�;�pƊ&�~d�9����c�I�LG�H:��K�����Ц+�R~h>
 �[q�s���4�^O���Q��q���6��45+]��[	q��8/5y�56���`j:���X������iS jI�#�q�"�ιjf�$V,��$ϙG"�K,��&�6�{9*;�'ޛ��G�+K=�'N�����R�,�\́3E����~�.�P����?}G~4���PBcv$	qd ��u�Ғ��,{�Y���X1���O�,t�_t�q��cl���Lom�6.��&�(�������`�r���ݎ�p��z�x:��i/ ޒ��	�R�0�#��7�^p��#��;#�,�G�9����rP=��U��?a���I�Տ�1}T���3G�ã���� P��X���%�M��}�{GFyo~���L�� �V�j��$,���C��o�u�75%�\��,���X�Wx1_^@��x>�=h�ʎ7��=����dު���>�ON���D���˭e�ƪOQ`�����oD�s�C�뱯ٲ[���L*�'ږPV���w� F@� ����:N���ɂ������2|n�n��Bÿ�$/}�ݫ��4�4�^�_��mI�iAbK+�����ʋ�<�X�b�������:��v�ݖ�ʄ���I���ؿ߃���}
�Ϻ?'���
�P�wW�gdxBt\��,8J��-pp���
����\��3��d-�8:}&!�����+���gT�� �;�nŷ\$��]ᖗ�T����C%�����%Y�
��ȗ?�Y��*�P��O�iI��C�	�(<�x�՗|M�ۀ�?�1�h�$7����G�=J�n�f��:EW���w�U)�S�Ի�\ɛ�b�>���_�@���R�_��6�R��u����d�KNֱ3v�2�xv��U�=jq�#�(=`�9s"�!i��gW�H7�9��i'�j0���� �mm,7�S4�G��$6:�WJ���y���$ sb5�^�)#�f��¼D.�`4�D��C�f'�c��|9�{������a�A֕p�缫G;�!N#�Cʴ[����wS�^v���)��ԨT=s8�	����E�"�
���G_�M�;��(z��.��gv��R]������%|Z�ì�X4�#p#p(΄�C��V��p�;�܃�Y���: o�ʪ��y(B��)=�?�e
�eTJ>o(m�[�h�1T@��&��g�*=��������u�)T���O�OP�w�4��"�V�I�XF:L//j��hL�����S��ז��o�95�v����1#1R���@2ɫ�@I��#�{f�Š��-��O�#��	,��{8Β��0����h�+�;�����f֨��[Fj�Ce2��Χ/K̀���{a߈��2Wע���1����pړ��sB���1�����5�X<p�F�������ҐG�&AYçC	��'�j�|���R/f���	Er~�~t�@�1�?%�y�w� x�V�p�����g����uQ�h�����&�xWw��O+��C0~�gX��b�����<C���َ�`�ֶ%�B���s�k�zi�q�-~!��[;�-1����@��~��_�<Ҋh�RK*Ku<�x�K��c)�I<e�Q�v[p��gN��ro�ҫ�[RD�t��Ժ�B��|ˀ�b=�aUJ.M3�"�SV�)�փ�`$D���{)��M�C79�W;o,�r��#�����
�����=�sM�Ӳ�s]���{z�~/b\nn.��0BE4��s� ����?HV�ϦɈ�k�F
��PQ�����٩WqD̹�֟ݎj�oQ'O�6�Q�E�R�۪�TD���ϠV�ƹ��M�C�<��h���ExA+����1p}7_R�K���a�3�F��5c�C�:�\��Y��L����Plڙ��M���n�Pa&VB��QV��k
Xk�J��3ð�l��%T����%��!��n���v�]K�9�M:��ό�uM�V$y	�q�}i�[,���;��
6�L��q��g��o��76�N�L�a�HkQ�W�C����s��tx���^J��R�n���7��cy����5u��VRO*���c"ra:�2>:#�[�Ȩ�nU��D�����+���7-��{F�|̯Y7W!�6x�3D�O��ʯ崼f���n��f�c� "+��`	w�@����ּ3p�B��4)�Mޓ�T�p��C����曨�٢R�*�!3��6�`�q��T��n��t�E�u����M0�O�[�^���5��:�I�@�������xWyw~��$�/@�y��_uB�~Z:G,����� �V��[#�;�j��6�� J)�߭H���ۓ*5��|s�O
H&%n�]E㏿V�O�ЛJh���+*j��<�Z��G?�g�5�X��������#���^yZ�K��o¼�7��&�u�Ж=0Y��5Dfyp��wHt��@Sc�RO� t����T@q{T	,j<�N��������)(U������Ě]/u'�!��f���v/=�8�z}	q��j
�n���f+�z�� �|M*V!�z�[�0�)p�֒�;�#���&QC�P�-b�Z��3�.������K�D,l�f�d4���SW��¢Nέ��? Wf�m��7��M�n!�ӛK��Z#j���y������h����;����ᕦ��\,����U�
���L9哔%�)�"�K��-�V�t�HN�o`���R�bҋ3h4yV�ľ�5��$�\X=�j�t��Jo0�{���G�#��Jb����G�}�!d��R5�bℲ�˄8�@���k�֏t|��p����Tjf��i��$R��	���z�����0��4y~��ox��Sl7ML���l�2;@�+oY�1CD��{k���QD�c�{ ��ϪFk6���,[U�J�K��6wWSR���Ѽ��h���$������bH'M��:}���'��tfg ���tS�Cu�Ӱ��9(�=��0�khB����@���찖�>ar�<��0�  \F�ݎ7�~ګ@��ipa��t�6zud�png���`6)1�ܻE9:���il�R?h�ܜ5��i3V��IJ<+ b �p��Ӂt�o2Bz��o�@��@������aA��>u)��"H�Z�{�&/P� biw,*�ϙ�[ۓ��de����^����U��<(�A��#tȸꂵ�ɷ���غ� ??w�7<Ml�HM{r�j���¥YbܥB��z��Cl%7���nũ� ���@w��e��V�r]��\_���㴤:��LKR}3b8���߉@�N��TҶ� ���y#z�Ii5��n�'#X9���O���tIo�����/�ׂ�_yhm�����L���ur�V��kE�-	�^3ΎJ��H���	6��D�@�B\>�}��rdoz�RH�u���*T`eE�#+����x����ͯ��_�L��}���д�Kh -��$���A�~��?<V�C�n�-��BRǩ��~6�l�v,c������a���j�s�N��4���_}-����t�6��KH�]�� %�tII�%T�"d3?����)|ޭ�Sզ���>���
$F5��jiM�\&L�A�_a}"�I0;�e�Mq��mS�C9z���h�(}�22c�܌Q4ù<P&JXX���b����<9"��!K�^�� ��P����d6��u�����lsC��oS�j�y1�U��z��m�p���o=���9~�����߸�g�5O��Vť^�"�����|9H�;H�7�XZ)������#:��JC�4W@�m�r�ܧJKڕm>V�"��:fg1|�K
���L;�	&n������c1�_9c-y
�t4c�)2�;�Q�v ����<#Cx���[Yc�,�0@ S^�9�4��Ь10Q�dRWi&=�G�s,mC�;~ C|?-� �Bae�4~�e[��{jP�d���G*�����:�+ch�r�@�ۈ/�Q1�5������)���M: �&���t$1���F;]'=AlH@p�g��VPΝՒ�B]���^���	H�����C�Y☁���b��I"�u���3�FV�\�ӫ��Yf��|�_6�@5=�c�mK��y]�� �a(���i���v��C�ZژS���y����{1�q| =�ۇ�;�S[���&��)���h���v���7��9�{z:[!��	��>n���	�H�&}��ӊ^�YB�G5ɸH	!�!��c������㵳6J�g�l]ԣ���U���8#q�/f��?Dg	 ?�o8E�T�/��	 �HZ�O�ɝV~|g@j�R����Y�H_!X�:pl�m��(ă����i���<�/���X='ӯ�����m�*���wD����
��157R |�0ԕ#����l���΄c�ntb�`�ƃ�}I������%:��v#�����"�>q�Z�p��)z;c�����Қ��\H
y3�Ѷnq����/B$�*ϸ�q�"�9V�����V�~U�͇�Fא�G>��#oD*ꄩ/!�-B�����+�<ǔ�y>��BN3�}�h�J
�KG`��X�ٴ(r�cZ�t%/,�=[lmRF{�^S̃}t�h��{�sS(V
���)�KI�?^���(���1"�~�DHrԝ��1�VT݂���8�R2���$�x\ڛe�������k�7i3����Խ��o ��ᡘ?��CRt����w����Ϲ���s-�� �������Ɇ�8�]�:Ƶj�����i��G��@�.����fv<��W�^ͻ�;�6�������|��)/O�\���%�(��	�����G���l �,�G�縺�Rb�5@_�N�a&�6E6��Eh�6֪f&��[`W�5w���]��䄖	�|���5yIԫ���S��W6o��q��}4�N���_j�3���A		�9�	�����'9�Ss�E�A���H��>B��+�E�#���j7:5��3��t����ά;)1=�+��,!�ϥZ��C㒃�f$��\s2�E� v;ID�;Q(�&v� �3T2l�x@��Um����aA���m�����bt(�hK��.�y@���D-��s��Y�#>��ő�`�U����I$�e9��O�0ծ�ɧ�ĳ�7����Cʱe#x����ڽ6Z�Ρշ�:��R�Y��{�A[�*KD��c�'6Η ^�}��PT�aG���㏣��T�IC�vk�W,�0�at�-r���	|���
���Z"
�Mg]AK �U(S�f��wXI�)����� � ����b������&�a��\�ȉ���A����џ^ځe��[��=&��w5Bw�:��H�$���DSg~[��G���t�F�=0�t��L�ϛr�}H�=a:��=�Lm�N͘�tT"�i4�Ӯ4��E��&B�kM�������,<zZ���$��Y�Cd����>���T���q�V���'�,�ƣ'�x�=�Y�!3/]���)Uhށ�`ن_&hT9��?�����h�����#f�P��k��$^���r��7������Mׄ#�z-�Y �hf3ԫ3i��̹��'�V���oeӌ��]��0l�M��#����I�49�r��z�
^7v5���͋��_JO):aJ��3xo��[}
R�?�X�c���ꤼe�%�wƀ�)��B~<�>�>I��gf��c����1�����*��ٔ�0�Е����T�KI�.��m��K��m],����,x%9Ք�=�P,�4W K�[�(�IF���;���m��W�=1�����7��������'F<�k|C��"�n;Էv�d9���_��h�P�Q㕒b� 
Sw |��e�/������{��p���T7�J�f�c	�ƥW�|4Y��|h����f|�1�=+��4j
ᨱXl�`j[��([���������t.�!�w���J9�(�:h��:a�FI���^d���3��e9��<0�g�Ӆ�ܖ?X�2�Hi��Ʈ����Mg��i�G����ݳ�X�'M�o�D�ؚj��=_	�;;�g������$$Q�% ��]&�j�t���P��}Kΰ��q�J
j�D�s4̪��c�(���
?H������G�L��ؘ�0�g ���gib��m��	��j�^G����t�Y�X��&���m�WΉCDK.����Ƭ@���T���f#q��������v�U��YZ����W���Ll ��俥Q�߅f�ZR���6�ePc�Z����Bt��pA[d��_t&�\�V�Pa��	@��� b�q2����k��_��u6��Eɠ#٭F��Pg�{�����YZ���5��\��� �)a�\�9:yk�y#˺�W/�w�5���7���
"԰���g�lҿ�r2/�b���u��SS�����Q0[N�D}Z��kJgA?�Wj� `��N�0r}�V�y4��f��� G�w
)(`K@�)�f13��WWT6N��xc]�b��Չ����BA���J̥�-���=����;�MCL�ks�%���y\�
q�*-/���� G��RI��b$�x�*��ζ�}�kbou:uo�q�C���/�]�I(;��gB����N(�����c*��"
5L�&-��c�~��������XI��`�jc���j�e�F�,c�Ve��!01�ED���7���'f���N�f�y/�W)�NHnq�Y`�ᤴ�>gְ��
'�W`��Q��%�i�;n�F)���,�A� ]���h��@e��*Jo��%��$�g3�i�>`u~M�Z�jz���Q��f	��Ͱ�e�Ĳ���hb���D��]�j����h�k���u�OlȖ�E����)7"�Q���N$b�6���4R��t�> �?�s��^� 2R'96�.=.Sk���%}��G�z	U��|;�|��D�rl�O'���Y؊jG�ն�^�T5�7�%xM�6�oeb�/�!F*\��Q�~��v��C{դqm�
c,? Ʒ�wOg�N���VL�9!0r�"��~�]����7uu#��-"(6��� �nu��iǪn���C�0�2c2���L1Q��ϽcQ1��]�ĳ�����u49}!VH��0�� ʎI�ſ��J�bf{|[*�I8A*!��ɞ3�w��<4C��C��ל�{n��/3N�N�2ۨ�qݱ���Ƴ��l�[f�	��k�0	�}k6��N���*!��d��	��C��Ѐ̿��F_)����&�4�`�@���q9e"?�ABλ�8nU��z
N�Y���옪��c1���~t�enߥ�-��L���/Vy4j -�e�d�a�������99awКٍ1����Y�J�/hQ`�,5��#����ӯ���ߘ8�uW�-�[W�㐡�����e�U��pv}���w��K�"���:����gб��^/~9��y1=Z�;l��hq_��l�����a��'��t�:�U�4��o��W���NR�o	I�3`��	�Wl}�Ǉ*�����*���X���x"����Iv`��dW
qH=�op�KI�/�#��0@_F�%��2��x6!0��#ϲ�Y�KԳv�v��A2�r�`��9U�=9�:�&仭ʷ0vڂE��e�*�"���8��,O!��{_оU+�ܞ�!�	0۸.�H��������`��MoOHwO1�?�r��+�Gh������ؕG���̈́u
�����Nߕ^g���*��OQ��'y�*F�6C~6z��n!�!���?�8�=B�Z�#KqEM\�$�܁5{NRϘyW<���#>�%-A�2<��D1<��P�1]���x}�՛�|&�zWr���e�����-��c\f�z�j��}��! Zh��ka#g�!Pz�[ ��<��\�C��!���M�,�%����˹��Ν��+��t�3���S��c�[�x�~�������rR���5�28h�\ׯ&�g�c�ͱ�E}���9�����Ԓ��"b2�#�n�	
DC
ށ��~!��!<y�xH�"��̤G�{4��v�p�q����t[�{�Q>en�Y�f�^��f��9�Q����Jv�CXe�)�DpZ���Vr%+F��w� ��@������Y��/�����A���	�_�W}��a�?|�)�.8K�j�/��p�,��c�Z�9�r|���[	��������U+8�ƨ�c �3zbb<��9w��K7���Bx힤�"���"��^�p��l{P��1=��d&i��u]ǭ�>�G��s ��$�s���3�}���H�v]$���	����Ӕ�=Ȅ� 475}�4�f�^����KNu�:�c�2G�wdF�����>�V���>4*=��Q$O)�?�o�������* ِ���7�LYP����z�J�	�W������7�n��?�):�~������<4h��WY��R�.k��_2aT,����ɢLJ��ox�b��樺n���.�~��9���h�HB��?�?��y�	5
���Px����pKq�+��:�:Wy³���-e�Q�_�ug�˗�;�8D�5hSU���ʹ�(��	X�'���_��E��s2'O��H�g���y���@J���R������� ۺ�;c���}ho�h��� �ۮ���5�f�K���������V���7�����Q��S�	�%��K�am�L���e��9�t�a�9o"�����1+��8$��\L#�Z��Á�
��֣���]qv�����@��#od{��*�]T��yJ[���W|6چ�'��V�e���ǢkOm��zo[`��V?�%Ȁ�]�G��O-��@��,\�Qe��_��UP�:&�靳�ħp�׃qg?�϶ר�HR-�x�劲�"Ǣ��#T�*��]� u�W���B*P퓦�"��S��w c�qM����ez����4��(���[$�����Z�B�v��\C�z]���C��k�����-�I�s萱O�Y�5�	#@�*�/�i-[�YP�Jjb��8병'������_g���Ay�C�[��%�=c|���H��1f�z��F;�)z�h���,a��	l�4�]F\��n"Z���6���44�W�`�^�cf�2`�B�+.v�C��y7�	�	Cf��5 e�<��`Kh�G��I�=U�y�&Bd��
�)�[^p4f�U���S7�P��%3�	�3/a�;�Hڶ�����'�e<�IoPh��lk�`�Cc솼��/d7Ւ�+��� �M��,�8��,��Iޛ���e��b�Q���Z[����m��8}����gaڹ���EpkBC�`O@n�$�2�6��[{7ԓŀ�8���=0p��w���h96��e�#gw���Iز�Ѣ����,���
M%ĺ�G����<^⇁�Ò�e����	B�"�s�x#e"��e�滆�D.d�)��:�۾-����C�ON���w��rȬ��W9P�̑Ce�������M�-71��]��B+D��76F��C���jcc����ZS�O���Sc9^�f�V���K
�v@6��t)���
�[S�}�9��V;�^j��7�������=�|�Kv~@I�ظk�^��X0��r, l��C�(`XJO�����q$7�=�A/�!���m�g���?�b�,�\8:���	��P�Ο�\��#��Mz��6o�Å+uL�#X{h�1. 0����,ʆ��r��9���h�kt2�K�+ӷ�dO�-/��j���>;*�_R�4����Sr�2F�5�X��@U����Y��I[����������?ϸp�\n��hW��i��w&�d���f��q��X�d�H.��򗫖���>��i-��N
�V��I8y!�緇 ��qĻֲ�K�t,�o#�3��cLQ3HU?2̆�p�aD�O��N�[F� o��������QP�&w���҃<�0ِ�޷;�6�I��j�ӆ���C���4��x����Q]!�'5���=v�k���P����RA�x*.tjS�����_�5�|7
��*���
����Jg��؞��3E"�\8��4~�HX���f1g(}d�U��jrG���I�-��JyO�jD��2o�3�2p@ !.b��M�'\��g6��2?;0>�\^����,N�fb�S���D?��FX!2$�.V�������ѹ��+<��aQ���g<P�V��\#�L�]J⸍gk�\tJh��E/��͉{��S��H*c&�����%�WH ��$��(�&������X'���:A+8��]m4����v�ۥ<#����Ԡ���` ʩ�@{ϗ�:a���ld+�^��t7�����(j��x�q�'b-���u1�/�*�K�X�r|(�)?��t�$qVl=��y9 d[�y�"�������S�m�����(4�M����"&̤��O������U4���C�U��*5 �G8�&��r�y���l����(V�8�^DIȵ
�0/Sb�a�e�.�т��[���8�*߽�M�X�!�/GR�Zy+�шھ���=�޾��d��.TIY��Hd7o/]���ү�O�a(�u�a�������x�쾧��m�0�4U����h�?�IP�U�6�͐o�N�������m}t�?^�L�ҩ�9�Tt=Z�d������~��s��*�I��o���Q���~_L���F[ 9���p�>��3T0ӱf�&�[�o���9�a(�N��7+/'�(Y�_�N���tRv�	���Q����ȨG�>�G�R���j?A�@'����"}y�fb��U��� ��S�"p�P<E�Ğ�8���Ms&���!�0��(��\4,�E����%WȪ����^7^�3��ؐHJ�e�����.������ '�3ȷuw�TKH*P���)!����~?�Ǥ�9����k�Ӭ�X�@"��|�| ��^]�q8��K/&+Em$p�"CG9�E_.`�pىE�Q���Ty�Mb��+8S��+`�>F��`<{�t%��?��d�X|�r1�6��A8���&��3����0���"-����'��	tzZ�f�o�ZlP��5a/>C�h�K�8�`N��gj^g��>����*�ٛƙq0�a{�ѰxH�B��dL�*z�{�����?��yē 2+����y��P�H�,�����ױ��{l"��Q��.1�\��w�9�ֶ"��g5�7s���E)�WǆP7/�{9���+���D���xa�H�|UT!M,��D)Seok�`�u���Lq�;�8/�+b�@h�~�/i�/��Y�hm�Zؔh�3�R�<�p�\'�p�8�<Z,-�3�?1�*���a?=MK��-+qxmY�x�y-C��e^*Y���nJ(�'�u+�M-é�S}�a���3�?�=��Qĩ-�+aaVd���-�Y��7s%B�@�ڄ�d�ӝPs�����3�)����a�"�}!a��e�������뀆)�*͔��9����:>{pC����=�_�;����O��(i��j��zu���g��̋�OF R.tek�æܨ�ʆ�v����)B���@���i���I�8w�IB��4�!��qm��ꠏ
�`QA�__��JR��b�.?�"�U������I��IeE�f�[�pk��Ǽ��夓+�x����?�a���Jɵ�~���%��)M��6X��HG��¥jMd�zaZ�^'�L����s��3p��#�s���d��$���bc5��K`�<�!)����6�3�|h�D�E z��O�2��~����.̸��ݴ)X\���1��"t���8��b��	q.~v�YC���T>�qrZ�-D�%� ��a�����ĭ~����tQ�09C����G��	�MkG�<R#n+��Q[���2{>�O|�bS�fY�� q�ζ6b���P	��f��Rt�t�/.��)|WA�7���-ͫ��k�"�I�C�v0����D�O<� �cPS�gWl�]�9)�ߏ�#��tW��6���Tu2=rC��9�|��#�m���%$��nL6ε�4S�ծ��R�Ht��k�D'6V:ɪ����f�T-���u�9<��nI�UC<���`�I�]��t�"��M=Ǩ,:-�h_ؚ8�%��Q������xƦ���Vw{����82A��%;^H�#s/�o�)���Ƅӻ�ǟ�癷I4��ֶ.tPE=��-0Bk�����8VDӿ�����(��J���5Y����]�PxJǾ�Y�Z�A�&P�}%
<V�����P��07�C8I�u\{N�{ ��EY�=������t�BL��mҨ�L����:n�������7Һa�ګ&�:7G�f�с���"k����,! ;�B�h7�5̥��_f0_5�xw�%niE���Pk/2r�l��`��/�װ���$R4�ۺ�i:ձ!mgwB)]ǅn��kޗ��Wμfb̫����o��O�u�_);>��j�r`"��=�'�nT3W�
��Jm�Y���,��2|�)���'P<��ZrT�j�ĸ��5�j��IPM*��]�YQ����L"1ɍ�y-���k��ً�4L�)/`�A���CoT���uj�$y>�_;�܆�9���55]U�A�� ���>bv�9��>	��	��7s�h=e�q�TOޒ�K���{��k�3(���K����Ȁ�6q�:� P<\�������IQlNyRj���9n�����i�	�UK~���p07W�% Z�S�����	� ��՜�/��]���TD��;q"�7�sfܩ=�)�qy3p�M��y'�%3zz޴��j�7�~H*ۓ^舁GJ�aA�V�� ���'�Ŗ�P�4%�Z��lJ�o�&�h�W����= ǃ�R�U5��W�<d�:|����b�t�����w�}2�攋.8tZ��,�D�\�*��ݠl��i�w� lP�����l����JW�AzG���Cd1��b�Q,?_�v
��sQ����y��e��T+�[gNy���Y2� ��U���������驰,-�OR������[�G[�ݚ5d�^�^}�t�y_+$��'b�+��r�I��0ց?c��ħ��#������`�!�o��g��N4 ��8w35�^(Xo'��,��\�z�XSM���o�ƸR\�2_���H���3��n�	�!�M��TY*ԔD6Z���"�	�l�������ڜ�>H0����l��$�c�3T�	���2�<�42\������ZܯU/�6bi�CC��"�KY�)DCt�:0�5�Q����
���|qz�H����/�񱓾�<�r��N.�эq�U�j��G��!/F�����G���z"����j3V�c��V���fYK�}���B���'���Ͽi3�����he�-�D����>��5y�~o>��U��%F�)Fɀ����r�d��L�h�6��j�:q��g��P�1(�=�4U �E�f������6z��M�(����dLOw�E����O�υ#_��KOSp,�����,6��)�DH_(�>c&�+Q�7%� >�}�l"m�1O���N��DOwc<��Z{����dx�������Ί�!��c�D�E�LUL�(�=�r��٫;�$~��{M��K݋m��kϤ���)��/j�g�k�73��*,�P�n#T�$F�T�l��	�"pܸ���<Y 
�n.A�ę�)�5�Ta.;1��,��04����ez��K9s�b�B�N*�h^æ��E�Hu��&"X��l,l�j�^΍s�0�ɜ�{��i�G#���u,d����#N����Ҧ<��~xD���j*�8�Ǣ����GЏ�܃�]��-9D��@N��FB�kl����7�,�]�e2�Yt�ޝڄ͓wTq��B���ed�7����f���"WnvH����
9x1���T��΀Q�V�<�)Z��
z�3Dj� �����3p����D�pY��.�V�6],�s�����t��l��ztcZA�1�����Q�h-~_�҆$W��|9+W~��'4��h�*�xK�m�2���&����c<�Ѥ��p�A����J-��;:!�
z�N_���~|�G��:j =_��$A���<?�@o���;l��k��,�I���m�i9ɋ�.���8���	fF�\�):�~c��"%b׬ܥ����PC;n�'	v��{<�,sj��ݣ��G�s�Ҋq.��O٭2<���_3^<!"@��pee��)D�R�7��% #�Jk���ob��Y���(V�=,����J�ݜ� �Z+҅?��s8&%Mg.�X0�:�Y�8��_GG��㺥`x!^�w{������<\tnl�����<Os.��15�=�<�	s�l�
/T��c��&�;����̒eY�&m4saj�,;�-�.V��cc��-�^Y�ϟ�QG��k�_f+�x-�P�w��%}4�����R����*֫�PBʳ/_�N��J$�n��tA[�����7q@O
%��&���!�a�?�*�?\����Dc��S��!Hz�J9��a�U���_*V�b-Q����/���4��'�n���Q.��4? ���iCy�8��������F
�+-f�e2�"��z�t?����diȃf=�8I��T�?����y<������P���3R̽C+tUD�%CK9��md�o���ke��)�^	��G���/Z�G�a�[N���U���n����j����9�Ҟ����wd�*ǒ�B�i�&�F�7�{�@�s0�X�AzT��L²�#�n���U���&��LE�2E� ���������ͩ��0��Η�%���畎��]�3J�Eb�T��r����H5��9㮵V��<��c�ʰ\�X�.5�� R�}&���������y�%�M�1�kup���q�u"���3Xd��=��aiz��v�x�6.��1	�]�7��ď��;��o��X�pRS���0��	'���>pHy+<�nЧ�o�huWճ��˟��2��]�Q k>T7N��A
�b��2�R����V0wc�#M���"ԗ3����B`j���MC�Q49���\���)ɉ��I�i��9�ji��|�]�|pj���u�J�#F�X��do�ʢ�z�
�*��D���+1�;i��%/fԱ�K2DΒ��ۀ	ל9Ś��}����|�^4��\��Oҡ��~�1--��W�bO�0�r�/��>]��%^/�o"��"��F��r����C`���7��[��:����nyRVkؕB�g>�!��8���SpɰE_�[v���1HZ��r��N)�[d/��A�����A���R)���z_��)�nt�f	�f��>��?co2������C�5��ϗ�6�(�IQ�Op`�V�I�m�o+;r�����x�H=���3㿐�oc��y���1HyF���6����m
�z��%f{V�Yx����`&{V�/U��c2�j�e>�b�J	�"�U?''��C�H�{�G����N-������&3��@��0�Ԡs
������G�*�Qˉ��P����ȻjD�O'	�&!vqp\�0���\Y`�t ^�(�~��%�Y���k�6��.�<�Y�JC���/�Z��FQ|o)˷� ��O��4R��F�-�e��T[!}Z1MeGjG䃯��b�1�2I�<�jQ�cDCJ�Xs�Q^�������K��ԉ:c�F��F(��Ʉ�J��[���eǲ���K7h�B���k��;�KG�ݫ�SUw.6�\r��p�
����S����#���L�L�$PX2��&���j���K?���:��-���da?Ρ_N����l��Y�c�Ł�<���d.�4�a�+�GG��-E>�y���;d����0���MJPͩ�F;��^��?�b�ɿ��v嬕\�݌�QA"P@y �uFXE��2�n�d��B�g�6�ث����S'�	-�a�D,����Kڲz�n=�@ܢj�O������F4��w�̱��n�اX��iDt�,�غ���(4S�]�)���C��6�p�jE�z���A��Y��^{7]a/V/��4�1Q�B(d� ���'��!p�~���,�E�hXT̵K�B�L����#��Y�{_����;LԆE�@ɯ�U6O*\�d��<}��#��F�Hr��8���T�va���&w�H����F���e�	���M͋J�.!x�]0�Z���v/����Ի��#���0V�����2�|0]�>�d9�0!:���{,�!��>��ħ�hJ���H{�(X{zS�!��y��Wz�[ՙ�5n��Y��z��h��� ��^��ـ�RY�>��f�K,�*j$
J�IJ0�a�&aOFc�aY�����1�zu��f�&�\��E���+��0݀�rePW�qz��u���_z�a�C�� ��D���B���˂��*nf$�v毴�݁��~_�\��q�$Y�{=|��(����ly��](P�.�������[:<�\-�?x�Ϡ�J�1r�q��N��=�n�G��OZ׼Z��A���,��%@����-�ٺnζ'�5�sX-@��c��&�^�A>D��I_��f�)���j���$���6P��\Vs>��SQ��¹E�O	��{fr��3���*�R�b�R�n���9�q�[#����a�kh������T����|��1��S�E8S<���/����㍺�*����:P�5&5�nPq�E��#��76ɫ=%��-�%~�s�̏U���G(�IyfL�pGJPѭ��业�j����q"UÆ��Bݒ�ֈ<��� �hk�ѽ���MF�A`X�s���%5Z���.��p�4�Uv�U#�t��=�im�<rA�<�R��h�Q��xD#�2�A!�+�L�O���*��be�`.�Mω$������(7�V�Ô?^��Ov��7Z���ݷ�l.q��|JV9=��FD���J�jpi�;tl`�3V���J��*��?��	.ņib�tB[	���ݜ�{�}��G8l�l{��0	�U�L�/�X4s�naAɳ) R#�=�����ْ s�C�nqx���)��� ��-%
�)��@�B�1/E�;$�(ף�=�(���k�Ĉ�LH�3�&��ޭ��&���*��Jݲ���Q}�a�O����
17|W��M�T�U�`W��w(>�����n��ꁸ�师º@�"@6�/���o�HӢ0�0������y��#%!��e{�ŐP�q�"/X���֟�!�pXH1�\5}�'9Gn7H�
��jIXH���@�|�N6Om���&�9Tt-0{ŀc���:��mӆ��7�#�V�.��&�@OMq�ÌG��=�/�hE��y��m�;�zO� BX������*&�#�=��i	+��J;�E8��o��E�ǆ�߬C����=S�HbH��.�!P���h�bZ����2��Sl�ҫ����=7;��+�j|�R��%��P���}���eJ�f8�(uV�C߫�!W���j'�R"Yf������Q�fMY��T5% �h���ԁ���խp0��3��U��ro�� ��>|�Ǖ6�a[��p��x��@j��ZY�yP���}�z���z�f�O�鑀�d5`��\��Q�:V؟i�H���z|���j2�̌�w�H���s/,M�VB;��Z�I�ǇM�� t���L�:�QLq�|�exL�&��	J�;uJ+/>��7-���y^I��SA�3�`��l��k&f�C���!��k�?��b�JXH��1P�3sG����q������1D�~����������؃&]�nZ��'t)e��y�m�3M�t��S��D�75�$�a��Y��N ���E}Uq�0g\Jh��\[uz��w��i���t&W+�^�`�mM�����x���\�vV�O���
 �p%�t�TKz���YVd�@ț�3�[^�8��K	�6��&@b�b�E��g�W�0\�O2��?i�+eu9��XŤ@zq���p� �_�J����D���3�;�̶m�t��*/�F.�GO�����z��m���$5N4�43"��_�~��I���=j<�����C�4h�]%��e�ِ��$���%���C��.���tA#�o�fz�~���������Ɲ	�+�
��G��Ҋ"	A.O V���m�,I
uw������y�E���� 0(6[�־'[x�`�D-Tn\~�� �"�E�H^���<zC`��*��6K�.����Z7�CT��=�5�Ӊm���T:s��t�V��7������>�},&@�bE(��ե�� n���*P%�-�;!~�i@�`�J��
����;s�s��Q�.2;b.?F��3"��ϴ�J��
;���􈀓�	Ô��Q�����;@�ɉ����MV����^�(�~P��"oM�i!���?��Ԩm*w��0� �di�_�8V�D�@�8��#�u2��l���
B�k:j�(6��G�k5�����jA9�wK�)�� S��h� g0�LF~Z����'�$�"Li +������Fd9��Y��
�^CUT1�ee������?�ҨO�oK}Y���0�viKwk�\�
s����<A�ѯ|�7Đ�lؠ%5)��Y�7"�ޜ�˂�D�3����R�?�up�C��4�T���zJm]�$����8��F$
PK��sGO�qdR�B{/q��Z�
�Ɛ$���O��U�ФB�x-�����pWN��B��XH;p�X뎊�;� ��c�PQ��u����
��iˮ?��"OV2�۽>Ҳ��b`�~^��O�_�����8�}�E�Ti(ۏ���3[,�PI��L�i9�D޾���F������k�ʏ���!a5��|���i.b�>��Iwt�B�C��t�dt���ʅ�N��C81h���4C:�hu�h"3�~�qt��P��7�M2��6y��sfT�I� �o�����)(���v'<%*�������2���[w�	���S��UQ��1�����[��6�~|1�g8���ԣ���v��j]�<�j�<奄z*ɋ�)�����{�I	W*w��F���&nGZk�	ǡ�ȩ��G{0JzN�$�(�:�l�6��ā��.�4�V��iQV���ą!
������R+c�
A�W|ؑ���EG�"�+]&(�xٰdh͟d�nH�-����ȯ[t�N{�ch������w��̖��w�Ս .�oV���%�-�G>r��2�y�������A��8��#���C��Fiq�κ;US��W�����Dn���T2H(ӷMb��268A��k�KuYq�4�3�|g�uė"��^�*5e�v]��pK?������5or��P�)0fl�X�lF1G�d��G񶘈O	���O�1|4��/�\$�ّ�ꍓ�Z��e��2�����H�m[N�(��4���uё�0�8� �?�(�:Ro�S�h�b�U�^� m��Kd��4߆�$��헅��hK�s�$vV��w?�il��£3kc�qgŃ��^e%y�H����H�2��U��>�0��; �A���#nV�mɍ��٤���s&�&�3��(b���%D)���;_����(\g}
l&�����Mи=�'R��Ȅ_�9}_i��-y+���?&�*�����m�-,@C5�Q��n�2�RH<��o���${�C�:r�1���lcUb9șf!���X�3��Z�.��/8�Ϗ+$��#��h��} �wI9$���$���q�Tm~��#�F��y�u"&X�.CA�Ì�]���D��'�ƙ5��_�:.|����Qt���y�=��~�/�D&��S�=s��w�ø�r��.��)N Ɂ�G���[7;�c���^��K2T:C^�4�� I����#��6�L�Xc������W1b��p�Y��xr�䗋�����	�Z�A�>���1�a�r�An�	���a�Ll�Gn���/���}Ώ��?��z2�����i��u���e=I�H�2� #;�Oms�&���%� ����.�|q�A<��K<ɹ�RW�Ǧ�z0�ZJ`;j[2�������:2�v���jc/�hD0��@�#�N��3t�MJ}庽�&#�	��̘��Re���<�W�V����]o���e0W`NBD����횅��ڋ���MA����.����5 /1��*��@�I�̾�n����,��;e��x&D����#����K�r{{8$/y��]AMd��z�a�>Z�fpI�_��r�nBM`#��K�񩱰���cw����]�M�?1ҟ��޲H�1�ñ���TP� K�v�ay�Q[_��HLkp\n�`b� �����K��%``�c��ͶC$Ar.T��
ˡ��~���8��§6O�:U�VzX�NG4� ����;h�Rc��Y 5�>4�+)d{���y�4t.�K�J�\�.�փ�1Qb_Ɲp�h
�lB\���Ԏ����;��nx�+�%�DW�Pt�8o�� �G&���ɾj:2U][�A�P\��SK�".��w�z5�]��}څ������IO���8�\� �OÇܙH���"��}��T��Q��?	������e�ȣ�ȯ<�PEfW��l��-.p��LO0�SɁD~�!��t#��ά�`�\���U_!�=΄��Z�Msa�`���3"�19^-Y�G���
�%����*�0����TCc1�;�ك>R���j}g�Qd.Kl�+bWl��-���9��`��H����������`���/F�v[t����'�~��īG�W� ݌>�o��ry�9+��ξg%m�u�a��E�ݜ:*7
�ܛ���ba8�l���������
�4;�ʄ���e��>�1���F�ϠAnk���g�Ϳ������1J�����`X�����uUf�!J^��U߇�A�+{_e�^�=>�p7����-I)����as߳�S*䎛w���;~�ƲZ���^S���-�+��?��/�z�1�*�)V8UpN����Ò�'����ܧkm�<�/�w���J�C.	~��GW���B���@jKUO|֓CUځO<������p�JQ�*l����p/c�� ��/�6���{��A�R�Ӂ,�Ҏk��l����bL$�۸q�0�M��`}�kz��v��!�T&�b�g�~�2T7Z������m/�Jɍ�����1H���e}��_�8l�岚-!8iԽ�
sM.�,�'��Xv�\��Kg��A�A�ں����yw���O��D����D�E�� 0�� �c5x�lC�M�� ��&.�,���*���E�$ٗ�¡I���>Ӣ��/��&��V �x�=�^EW2�y?���q9���ZmF�P,�7Z�O����d������� sj'�����0s��(7sn�J���u� �w��|U`nش�Ū�V��Ѩ�yJQ�(���9�]B����Bk���x�"�S�@�7���#�>nQ����m�������%�v���F���:�őVa�j��JY�_�'�dmw�%/j�Q{��P�o=���܈�Fd�D�<�?��uS�q�!^�?f�]P�' h}�����3�5M&� ��#�Tvn������j����7�F��Ug�*�A[���p��h��W"����#��˪�"�f���_�!≰ǐ�����i�)T�q�4=�=6tUc�!�KN�SF�t���ʉ��|��΍7.uD��oM6B�oX~�p���N*Q�&��ӹ��<�����P��@�/CMY��
j� 8� &o9�ں�f��{�¹���*����hAj����+��^������~��\����v��l0Q�[����]h�[�2n8�u^z�e2|3�}1���)��of��O����a!�d:ޖs�i�x�I��p(�RO�}%E����X{ �f.��PhbX���-�
-�Ę��e����wW��%Yt��lƢ�	]����`q�{{����=��ɜ�t�.0�f�m��j�$!6�3er�'��֡����.UP��Kw�&���7CLc�(�U�p���h�	�sZ.�K����� �垧�5��,��p��bR9[�k/�K�6��Hr�TM�#O0�la�8D�aՈ��.�pN�c�;���B�l�.ܹޝȁ�G�=:5��Nd�<ݒ�[�v)F+�$M�E~���x$}0Xn��L�;>Ij���Ѐ_/t�B���#�@IE�K��u1<*)hʳ�s��j�п�,# ��g>�@+�-�����n���U��f* ���x�Ỗ��Ac�]��O� C��Q�yB�^(�Zer�m�M+��Y���o`��*��c�c)�|��|��8���P�{�	��>�w#�玟a�J@��ˑɹ^.Rz()���Gf̏u��] A;��1r���u�-�ߚ�y-PY|�|2 ���� U�t����*$���՛��1C����;E�t��m��v�f"���e9��5�X�|��-��=е���[����h�D���[No�=���ԕ x&��􎟁r��i<c˛*l���2�v�i�!�rK�z4/��FR*��HX<����B&]�-]aK�������(���c���/�0s;��S�^���`����wArJ����"O���أ�ϻS9u�66� ���J
�V�L���4���M�gő�0�tȐ&8~/�i�W��: M�%&!t$ ��2����E�7Ҽ�g�<a���Tl��<��$E���Ύk�S��P����KZ�"�i��؀���G`�EC��n ��H�i'8E5�"�(:�?E��@�������dRi�oրɫH�0[��z�k�//��r���>\`S���\�|GV+�S[6�Ք���v��cI`�������;|]̄0����`Fh;�0פUr?�ʷZh|��[��ՒFDM�߽�5�۲w�j�[���� ����6��yI��Y�}���?����������p�W�l�����A~C�v���P��m��؞^Kj"�D��j_�k��K�у�G���"����wu�ؐ��6���������~9�z�x�Y�
��Z�ĩ��D�S�A$���� �H6��V?�=��N�m7s4��V�7�����v�(�l��c�;Y�.3�����
W�S�9��;
_�L����v���I*u=�,��y���\�A��ȺZx�[i�?���H?��;<�ka�SS�.9��g�p+�zQ8u���G����|P����#j�q(��,���_�#�I��mń7��ڜގ���+�:=�؅��f��f����	��]�9~�7��RPj�<?��d{����1�U�S�SY�v��ϵR��|���*!�d����}VΥ�~�]�1�f��w!t�
}����jM�H4�:m��
��!"�4CC�z�Tb��}S�D�
r�;�c�-��86q�F֍tJ�T��u4����2>&(�t�(^��"	�[��R�vq�2^�4�Z�2t5Ք�m��6�rvr���o�F>��ΑҌ��{s�<�j�9���S��i�|�=%�BIi8��cI���E|+�K���{2մ?ʨ��C='X���;�8��:m���lP�i��V�:Y:"){9����Q����8v��@��� ������Ɓi�FHJ�C���d"i'e�85��.����^�,:�\e��mA�7��Nh�
�W����F3�8Ȋk7�[a��A�X��;N����r,ҨZ9s�(��m�)�GWh�06|���g��zJ%%9=(�N�ƿ^b�'+1�gb2߬h̫i���a�c�X�;m�S��),O��_��Ut(�����򀋊�H����N"pVz��M�P~z��TM楉^��oX�@'=β:^�x9�|�Tq�5N�얌�K0�t�J�ș]� !��u�|��Q���Q�sk	������ׂ�W��9e��#|��qhr��}2x�L�c�ۏYi��;�S$4OJ8]�~��e���d�U2L�&��p�$y�tUg��w=ذ͓������n������@��\xN�w9>�e�g��P�����E��
��/v��W�/r�)��{a�+�QUW�n�2]����	�e"@N9M���? ��6/āʺZ[��6J#���Z� 7dQ��ks��-Ad���x��3 ���y���3=�iZq���8R�����J��%���^����z�����x{�q=��eeYg�P0���A��h��l0q�:%To�o?3�������(G?��^W/�\������gK2���R~(��ht;��i��'^!�B
%δ����+�敖�U���FVY遬jU-d���-�B|,�Jn�ɉU0556��=�^Jw����s��w���Ø��պ~ʱ�*�"hg�{��d�p^��o��t�ܓ����L�h_�eϷ��e��|���CC�(��DJ��R��RN�߿z�'t�M�h*�1H7�h�^�pz豀�Z�� �J�"�����ͧr��E��fiMjB�>t�=��u��i2~���`>eYw�b/��yd?�"�w�R�F'����pÐ�{٩ۄwU�Q�MO�κY�O�H�t�bb88���m����O��KwCs�b���i��|@?�����V=y��8����B��N���9��9�ޤ����ֈ��� h�BG��)e�->�j����N=g���=�K�/�)���잪��t�Y~��1�i��r�u�a�Ʀ�?pU��2鮙ԣ�@�e����e~��~j�'C��r3ax��hCpöE�)���"K�o�E{/�[x*��j ���?�v ���\lR�v�[ߩ�� O7���'~ 9z,u �U����"��C1~-��9�`���s�m�0 �$u�P7���K��R��j`��$r�L{�l��c�F���9�p �r#�������Ҟ��$˭#-�?�y��-�1gH��v��(n1N���D��`d�:Ԝ?����Z��D���NH����	����V]�HsO3�Δ�������$qM�Q�����Uӻ����>S��h��bF5��cct���D��uӷT��N����u�.|t�Ƀ�m� P�a�q�.~�&k�����ݻ ȑ�j �F�B�вX$�jk�N��,tb����R��F����ݹ
�k
���ø�L�6�q(��|�J��*\�]8�.m���Uo���Ҝx�r�,Բ�__�E�vׯ�����82� �g&j�_�%�׋%e,�j��Q\�J�S�����b'�j��y�5_|1r�6$5?*�CCm�,xK��2��a�=�\3�a��(�ş�#7�I@���w-�PaK �ʮ6ZH�;`�V#>�1�+=мV�D��K�*$��fF$Qقao$yCt�s7`�o ����<eί=�vu0�����&�Ф�:w��]�h����Fƹ;��6J��i��I�f�6�x��{���2h5I6Lq���Y�q�U(�ɼ��_,���`�2[_�G�P�����RX�A�A �1�-��$��5R>���x��`#ݹ�z����M;���`Q�{�G�X��ғ��s��o����蚝t�rX���6�(`�UT�f�d���l#d>~�i&	�0��5�/?b5=`�����pr������M7�puׄ1J���c�ٹ���I��V�[����[�gAfy�ӫ�L�	��vc]ĵ����0K^�?=�E]�Osv�DL��,�L؛���)�uo�z#��y����ĉ��gօ���r)�Oȥ+�Ty��+�R�b�ʡ[�KܩK�@A�Fzs�c8Qb\{�Z��k���xx��gk暤"�6Yzc4�f	��B.��J���R�����t�t6����Y�aT&n��rׂ���7�S��D�;}Gg�Kok�X��)@��A�Y��N�7���zw�O��4��@B[XC�7ip��J�H�F��c�F0�F���1Ed՜���0���r��sLT[4&�4_(�5Ο�՚�h�S�_3-�z<Q3t6du��ŽF��(�X�`����8F�7�	1�V�z�.��!���5^�ޔi�u�if^�>8��譵.P���B��9�쑦�(�3�9�+�6���#/GyL�sb�ȓ%/Ll|?l�8�)�]_��Qd��f����U�e��[d��3^�������L�3?���HE����ݔ��� �}���	����^k��	�{x�<ԕ�,>d�7�YJ�5������	�o�Z�βy�]�p5Xq���2��|.�A,���bC_�_���Rfι��x����H�[�S����77.�P������=hsqc�!�zp�d� ��	%��Xԧ�u9p   �R�C���i�Q��[����O���U��4�Wgs6�J���I���T ������9$�z�\��-}e�� aIvX>�'�{+-ڵ��s�O+f��%|��n�:�?���)�����9bPo.���h3�z���c���~����IW�	�5j��L�Ս����Y�' �q��X0�o�"��|���FS���s�����Dk`�����u]O����1(�ųsF�΃c�c��MX��;�a����� �1~����@+ w��3,Ug�㝙��J�َ�g[t���@cCD���,aN�l3|`���gWeN��'8�&
���S8������+D���=���%ļ}��Y��J��h�T;I�/5�H%�(�0���J�h$�1S髕7��tX+Z���̟!��.g�>�V3ŭ���U� !�k��}��G`�?؋K"�}��+�����8��t?�V��	��Y�nM_s��g�X�-�F��8���P�M�����L�
Q�����q��1��R�#	��@AR�/d�a��VC�c*ѥH���}8}e��|#B[�
h!�Y[��y--=z�p�Q�+?OX��V�UlS"Pt>�����eۙ�
�ք���t-�I����X��Ad[���u�fqZ`�*s��E{����k(e��{�,G���6<ᘪs���+�]�P=��5�3(鄂,r����Z���L|9;&5�u(�K���߯q��*�N�ߘ��[�����	��:�j�e�%_�?�:D4e��"�J�����u۬�^ǀR6�^�y� �o-�C�Ffd��F~gPΟ������t9��D1��|�@��C �D�		<����܈���T�.���ó�^Gm����fμ*�~��M��a2q�QEa��(�yG'���9fW���)� q!�J��֋'�z2Gڒ/ˈ$����vh�X?���v�[4:�v$Rv�0s壥x�L�N�[dn��4]�WsJ1vK�抒�5+O��ŏH�<�>���i���0>}�,?_�JrhV�y �a.V-����n�ج�e�A!T����SJ���su����1n��/�s���w\U�a� &(��୛�
��t�sS~�W�}���v��Pb���'��ѐ@-ۺb�9P�����LO�z���S�=���;���^lh,�޴�f`�aq\Ņ���nGZi�n�{Xth��!np-�H{&e���>��Ȓ|ak�����bH�9Zꌈ��$��~��n���A1��J�~PɪD0l�+�y���
�p�d�*��--]btN�:�h�~5��� A�U	 ��oD"��k���qY��$��t*��1>�5�v��L�#�);a�p�.^7�5,R
�K^0��:U��Q��nx��a߮ee
��V>[�t�B����Nh���ְ������h��n�̮ �u��:knj}�#�*�
��-�Y[u`n�\����l�6�YmDE��No�po��;{��V�.o{\/Q)�{3@�$�B�9��y5{{ue�V���%yfԚ�������Ǝ{ki��ll;]��ig�P�5$����E���"�3�a�[�X_������Q��ɐ��w���Z���b	~�8�(�/������υo��tl�!v��@�_�V�2�N�E�Z�{!9�p�	E!B��t�ӥ�Pn��
A7��ep��pX�(��~z ߱iu�ZVI��5F�]�i�'�����5�S�34#&���Bk�f�^��Ef�����b�*8��b�X�m�-b�n �>��R�A���pqe�����*��7�T���Q!�7H�:I�Bq/��~���RI�.��\���c_�����ʺ��Z(��*�s�xJV\�͗�y�!)�p�����B=k���UP�#O��b|.�@�f.����C��9Ueo�7r6�]���S1EE�������Z	N/}�p�$��
vqF�%|�Q�d�Qi+�w��^�ٱ�Z���vy�U+�<��DtdLG�<����w�^��9����iy޹cU8h�cY��rn+{��"�$^�BƜ�((�ꗮO*t���֒�����s�	�ُI��P�m�rW�2����4,�5C��𯭃�����h�;ݞ�g'��:X3|�z~=FH���>>��w	�-��=̃���?����5��*��*��R�7Y>�l�R����p�xMk��`D5���
6�-�m�ȟ=����v A�>���P�<��;���RP%�)��lH,��giJ
�ی�<D�dEZ!s��W��{����met�%��.N��̈Mk�_O&�M��[�Ӗ�䦇�纈n93\8�E��zb�GaJR�br��׸g�C �zAt�s�պ�OI6�ٛD��d���B�P+���R�8<G�ML7ʊ�L�AAz?Jt�_��vyc�S�<�e4�ќor3�G�N���@�N�|�#�/И�������,e��u� u�_���jP��{0�V}�,�j]e�ƨ����&�4��K5�$:̴��[�Ȓ$�7�u�#���qW�yR�a%��n�"w�@w��x���H��*_C���	�����%��Z:E�7��To���;a�J��a|�>�f��zgm�18)ۙ������
�/fU1�mHl�H�uej"Ciپ�5� �O}���!�L�'?[�*��D�N ��[�6�Y��g\��F�ܦ}�9�+jm��@�2+�	�F<_*$T۸�/d��/�m(�d��~�k����nf���Xo����]5����������j��ǒ�S
��?�x� ���F�ȝ��V�?���ϲU�;�6`W��71�yK��c�+�}ٻ9��*���JL-� SM��3���S�IK���Q�I��������e�E�D�E�%�dmx�����[RyV���~�񘃋;���ؒ�7��7b�gv��K/��k�@
�ߵ0xo�B��Z��+:���s���Ĵq�W�����\��j��ߓ�?t��Q�M Ui�p�@�Gz㍢��`2�ּ�8mo�;SB��X(G��k�#��h� "�+厖�Y>��xt˲;݄	^���P	����6و���b���g���	
����#��}�����m�� ��J�,����yGy^
���tj��(m��E
]|�'�2�4��&�p��$ĽZ��pT�B4�k�,g@�S�D�,o=�Sz�2ͫe�ve"&�?�@L3�l?�{�n��7��xI��i�����k<��>��e�0�S�9#T\9�K����39��Ovu�Ŧ�B�u(�(��o�*y*�c�)5y� �t�4V��{_~j��h�M�'��DM��h�a1H�79qlRU]��+ՙ�UjJ��bL�%0a0#��$V��	6C�MS�	,
K�X� ��(�+�)�)s&���w/L�i:����CmG��
&iW�Y$��1��D����nNX�$������<�:󫵔5��%�9Y�p9�[xk=K麏G�N�d��1+oс0L��,�~�cƱg#��g�\�X��bV� u�w�̗z#�����ձ>�C�4�jFQ�O�|| w���!���Օ��:���i8�E��C/�0r�H��)��e�nr|=,�v����j��6B�)��y*��=�eHF��L8j����h�X���K�m]�m�c�	sw���U��:���R&���l�\ZU)� �6��wOsΑL�!>��xL.�0�Z��7R�Z�2��L���Yx��m�r�1��^�ڔs*�%���S�M1���7�e��f��0��K�9�	Gpc"���,Rؽv��	���&�Dwvu$ǽ�FCf�Pb����XS8o��̞��u�a|`P�}�2�Ta��"���7�t&�:�lŏ#�=>�M�D�t�ѿ�v9qj25A"�{RR�a��;�tQV�@�#�=q#�v��&H��<��d/NTu���yO�F��Xvw��~,�A��ޅ����:xg �m=�"wz%��"��?�C@��ʵ��R[����_��D�Ð��7p���Qi�>y�')�
��-rH���96�슡ڞW���}ƌ�R��60f�%�W8p�s� �H�m ��abiĖ�#��5�W��ضJ���_�Z�Z�*�>�%���o�.d`	�����Ρ,��ܶ��M�����*ع��̓~&�j�%�?��؝��v��I���p�+�������άE(�1�����)Po�xu�:O��"06)���'�SB��w���K�W_�Ɗɋ�nO�|�t�	ѿ77��9?W�j�B�f���_�c{݅~��"�s��p��|�����BZ���٧�l�ѥee��#�\�: Q]%sqb�����x��J��פ,-����p�ߧ����?���O[�p�	�źd� ���kΟ�"$����(4g�I<��X2��Q����ܱ*�JMwڤGG�'��w�r .�h����!!�A&��&�󋳵�+ף���"��H�vk��Ѿp��i�]�9�����U�V'�B�S���M���I&'�
j�GɍR.��4�{�|���Z�k���Ůj���El�o�Npe����$W7Lb�;[�d�z��!�4���?0P(�uI
c��p3Q,w՘K6BP�h-M��F�H�>.硺M+g���XJ��v�1T̮����8�Ʌ�C?WH_l�u��Nf����g�K$/�(�1x�
Fi:ɶ��������{��ĜT]"�Bh$��/r��R�&��(�%v��3�d~���ܠ��0�n�̃���J}�y���`sa`ʏ��Ϊ�"��L!����*	�·B�s�ԙ�����A,�8/&o���^�YOC/�Y�.�����)j8v�|sE5�q,'&P��	���,4_�x��nٗ�<l���,Xp9�`%P@��I9fi�*'�$�j��{��N騮�Cq�>��`�G:?� �؄K[T��F_�v���Fw�Nd��r#��a=���s��y��6��Ѹ��R��d=v0Gl�+��/���y�Qg즦�͞�r��:�uq��W/�b�ʹ�Q��Db�H2����>=�H�x~�h4~:Uc�a@���ܜL0P ��8ad�{T���L)�~��X��1��N�N�5n0�V���!�b�-Y���);��p�R��R'=� �����!R�w���K�Rү���e[�EH�Й���걱)
��\�#�U���Z���}|o������r���ApTyW�w[!����nj5xs)�C�^�/;���<0D��!(�5}_+�LC2���ց3T��mt�^���)B�ɷS{�ǝt�DC'%���*ajff�r�0���
����z�O�e{���v��5	�����0��bǕ��}��:�vd��l�N��_jK,�Ͽ�fe��.�k�[���)�ܰy%A4���d������h�Cͬq/sH�����!&�m��O9~s�B�7�r3�^/�N���O�4�� �a�Q��QS�������!�[�i��y>XF6�	�A�k���F�X�u����[�[��9�:l�&9`{�ם���(�=teX�#t����8����H��La��cr:J*Lڤ`T�SP-.�{X��9#V'��7��h���?�?�>��$�r*˒h�	?�s�+���H�������K󯹢��k��"v$�zFO	3i4�U�I䙅��EKx����� |��xv�M���;h��"��n��&*H���'- DZ-�NytPkFW��c�P�1j�!V<s\�_p 'ܰ5�(��x@��Uv�u�1v�xR�2հQ��h�TU��"�S����V%@�U�͵YŤ����:�H��#����[iSm�����[0 A�[�}Zgʉ{����Ǽ6�U�r���x��4�ӝ��EOh�/�0n��(4L�`�/,�e�����w���'k������SL y#�ty��������S�Q?������N�m-�whf�t�D��&�G�� ��泯��;6�f�E�p>�Z݂G���;lF��v�Q0�P���ȡ"�,�m�g��ϧ�J/�0qvo�sU��`�0�zY������:��@����<R��H�tQ^�f��F��TX�G�x3��ޫn��)�ۨIZ`� ���}ފ�
V��xj&�|�%z��Q��Y|F��
�]W@�k
?�Em�3��n�fm�>�t��e{תEX$�hQ��E칛�0|G���e��_�sF:�#���,���>o�w�z��"����f$��hc�E�q&:�5�l5���F�rBnIТ�DF��ȔNB����I�o2��<ש�H�m��"�Gm!�壄\q!ւP����M�w*-
��%ώ��I���Yh�HtJ뭵ǼC<�O�"n%L��z|X�T���G�3�<:4G�dl҃�����ŚbQ���X�Xޚ�o��6��
��Uc���[�u�԰���'����©eg�Bɧ�~�e��`�
����-y��N�J*��>b�WR��/�s&������嬖�����2^��t!�6�:)��|�ރ�E���j��f�6̮K���PA(�95�͈iXz�����(�y?�����9����-l�}Qf1�T��@�Ei@�ܤ&Q
��O9�(���5h,�x8K5Eg�po#y̘��>%`Պw�u=����u,XY�����s:���=QY�̖�W����	��S�0^�V���@B��x5������?�&!�P�<�j�<J��(!,-�p���04���۪"�y��4���w
���t��N��Ro]R�0M$��̡��<VR�t6�Z ����QP�k�������S*\	.����`PX�=�LԆ��w͊I,�S�bA��%�63a>ep�H���7�}�bn{���c��G�& bژ1*�h|�.b�����,��L��j��<�}��"Ų��^�4��V�
o>�Y�����,22�𲃡a�s`�����]@ll��QS4S:���vU��V�$��|�[`�?������9�$,��'ף�$���2a���A= ���a�}���4Ǟ�)F8�IJq�e�	���)F!�FזB��>�33��ɡD:�0�%y��1�Ҳox���Ze��ƽ�vw9-F�KR�~�Ö~���*��%;�c��P���tO����:��7�8J�%���jTf�L0���8���*ڴ1"��B���F�G�b7��OL���{Wi� �@��RCV"#k���7-��G,6�4��i�����	�"lh�/�,��rx��_�u���s��dT�~�Ok���+��{���B���^D��|�}f�6�͋��r{�@`8?�7cx�_�2�b����������8{��6-��]-�[?0�B@��F�c��KTPTa� ��ݥh�r|'`��pŜ���BY	��U b�4�-�a4˹�����x:N^(H/�s����.�'����^MX9+�����t5U��K7-�_6�g�������,�������@�-c��X��ד�*ȂR쬠�k�����S�@����jtg�K0zd���`��j� ���:�a4M[�?���{H٤�:[��u*�el,0�j�6���6���kr��!����؊�&3JJq�bZI�R;��R����U�ˡt��ؗ5��A�/n�l�yc���R�J�Xگ�_Ux�ș�m8����e�1��4�@��� ���M�|E��k1��"�\d�����e.;��"���Qc�擔iWN�v4$Z��^~���)�=-݋�7�r���?Ī��,�o�v~�َg���t�şjU�����Z�7F���ϻ��^a٢��y��˒>��@v:P
T4��j!��9���A�ۖ�������t�xS��K1N@����4`�/s��u��32	�?疟�\�d-�Wm~;��
_�4�<>���z��եs�	l*Gd�|��cŭ��9QC�&Iym9��"����S�L�qyN*�ڭn-�����K?�(d��-�kB�H`DyB�Lǋ����1`IZ���v� �u:�B��5�o����h�'�܇hg�m=�;n�־]��d��>C p������//e*��90��GEue"8�M�T�4�X�Pzh���pn�w��'��y�B��J�D������v�!'!�Qe���p¸�r���\�f��)�ڔ=�^#��d��*�	��8
:��8\�Y�߁�SEM��8�B�n�n�������sIrZa�b��v��hBT�-�b�":C߾��H$5E��
��]�����i��\i�xw��+l�����3Y<�O��&�|�Q�-`�p�9L�x�f�LrK#U|���Ά��z2zݠI1��B����y��m+R���4�8W��TH����!�}T���`�҂����6��姖H�w�IQ����-�3��|����_L�3��_	~(�Tz�"��ft��uIXEr�����	���ή�8ީxr��nk�ѴZ�	��y�c~�ktI�����q{r!y�n��y��|u��r悡(��\��Q&�_6]k���ˀpNRv0�=q��:eR3��d��#B{|*�;���[��YV4�������q:�����0� H�~j�ry���԰ZH�*�/(�GNW��>� >k���N/5=�lv����o(���9l(=�.���8/@&����f5���f�D"�!���\>�ѡ�l���+ߤ/]P�u����	m�{L3�*�����Wm&|���xY�f�>%�a�^��� N�~%Q
����=����)6j�I^s3iP�!��
w���p�1�;ԁ�S��}ғ��'�|�v��MQ],y,B"'�_-����YM��7�.bY���2K�=d�(u�?��+�H.}�۟��� ����ƣ��~�x�g<UIP��$R{��V���*(+N16IǛ3#�x秊+׶B����9�23nӗ�5O��̾ CԜ�-,|�W�ᱝ����2f�c����\��py�E����787IJ�Fm�/�$�mE��\j>�c�w����9g��\k�R��d�W�#��:��}��$��[h�U�0q�4�b���C���I����Kdz��X���ocb]7/�GS�^J�}9@�v��L]���۪����j�+C�(��G�J�7�]��

b��TpV�DʦJ�_D��;2OoYޯ�H@�sQ��Qۻ��[*>��[q���҉2�W7'Y���N&.��::W���2>��k�#�\g,ã5�����u�����|�?�7~�����EC�d�և�UK��M�n�dJ	���[l�g��������1���EaxM�����)�r7�I���c	�����V#Y�46>�s��%�ڧRv�Lm��7|O��k��8��S>����3H�wI��4C�����Ձjr(��0�%w.�����%��,���c��N=���IJ��X~�^�\�Et��T�#totk�W�s�o�)�~�������C�wL����^����#��>b��4c��))�S��4��D�o֓~>s���Tȶ��pT׶��j��yVk�o�}�˩#��KN���12������v�:��������]j}/�8�N�}5�C��LÕgζ3-�u=�``U+�"�^�O��',��?~�N_3�
?l��*QM�����؀��g�Bp�y�`��+�C��5�b�����|<-�gD��6�~$wJ�}n���9��֐���.�!�sFC�oO��!4�D%@��r�������q���?U�P���ywD4~�]~�t�X����?X)�\��KCj菀�>�0fi��C��C��=�=�6�@YI���S��{�G��P�6�ӡSM#�[u��}&�x��=�Ĵ�쵹�a����*D-x��������|��Rƪf~:/}X��sH��-@)��p~�����1^��]�~�d��y K�S?J�Y�
<1U}ӓ���I#��܁�~;)$��%*v߉�N�<�������N���5�3��4���.ܵ�*��'��'��Ħ�䔪<쟑�a �T��;s�U:xI�
�,��8E}\n���t�G:��q/�T�-X{wEV_?�q�L�r��pX�v��i]'0\�*��D6ɀ4qDӃ^@h?�|`	?Gܵ�:Y|S^QNcđ��Q3��vG�7���cOƴ�A���D��_��e^�V{��bZ
)A�e�a���B�8؃}�i��x��ܜM6Q��E�C�}ȏB�7�c�q/`-�*���R�������2�* "<Z+��X>�cdk�@6���4��2��/�V�+28��W` ���T�vɳ#����A��d򡸐�Zxܶ�=��_��1{9H鶠�j��A�w��_'�9T,L:uE)����I���F\�"H�m�n\�D����z���Fd��GłB��J.�7��[-�GRƺ���KVnL|O��u��it���Ȉf�hE?��OԶ�FO�|��[���.�M��U6�2���xq]Ȗ�j㳋������Ġ"C�>����񫠵!R!������^|P1Sme�3�$~��J�ܣ��D]ށ>_�u1���3#��6Ƨ���H�뚌�h:ip�_z$����+7�����e_3.�|1A��z�2��>�qȿ�\.8΋h���V��qe�Ϯ�P���Ԭ��)2~���~.���&؋!u>���������F��IC?����~���~=���0ײ�;Sֲv��x�G?.2��Y9}��1�X�����&me�R\a�Y��1RO�G����U�a�zs���)I�7!��zԕg�ap&�u�������+K-�7���ɼ
m]��!�JH�Q���K��Þ�$RR��v}��q�\{@�!�-yԗ-�2t�R����P�n���3�-jO�=m_%�)���3^�s���b;WFϲ�.�Yo #�J��l�gjDR��xMP/�>bzZ��d��5h�E�?���}��Mp����RR�H����t�r�"��J��G�c�#+��b\v�� �D���K�E��_m�4t�tm���f��x#��U�b�'���>�ʃ�|Βf����o�RR$�*� � l��n�"G��Y���6���X�K�;��cH����jM���5���3qoa��c�� ���B����7��O�:e_$!����b�U�Yf�.?�Y� ���K|b�?�i��C���=��-
����).[���d��l�UR�Q���H��n�6���3�TP"��E��X#Ù�D ��S���]�: �����Kl0�����4����Ȓ:� ���{Q�ߊ�qڗ$#��٬�'ߋM͐��.1JMj�'A�� boȅ��a*����ӂ����}GE<�El{ Cх>�/|wHk�S��`�p�Q2�W	O����w0�`���M=��B����5�m[�C�aH_�����gp��7=h���zN�"��7R�7JW� n�p�ỳ�����
��X�#�����"F}B��	o�҈�x	5����@.���nJ�9d�Ô���K�kO/�ʯV��L'�?!t�F�L�)r�AN$ܬ/�i�L(���[�s�'�d���!��8(������ �x��%%;��Ǆ��c��9�t"�ŲZ\f�X�ZJ��� �Tz��TIcw[��<�;p��t��y�����R�t�"��4�K��9W��U��o����	T��2��Z�j;�q�>�:#���q��Ϊ��y���Z������Z?���c�HJ�2D���4��ꧬ�$������%�\إ�21���W�]~�vVW7ܻ���Գ����s׶����OrV��y6��ph���
4�� o�M�Xc;��æ\�5���i���P��Xtsg��
ό�D��E�oـ(�G^�˘EM�p��ս_����Z��圵3\�Ķ�DȻ�(M�Ͱ��}���2�˛�K�֚���U ��-Q$��ϚK�G�s�(eI%�6;k�P���bWi�\�g�M��i'�*��J,&�o������c�P|~v��}ҫO8�w8��ݲ�(N�VS,R�����%YL1^x:���?��cUH��8s��#�b�r�-�nf��V\by��a�YΪ..�E�\��t��ΪT�ꘄkw�[!5tfF�"��;�64]W�p����j7�%ʁ�`�DsWE����a)z���=íD�܂������_oRX_���x~^2C>u�+�6�#����tM1p�o��BU[Gs�$����o0�����,o�l�5sy���z�("%/v�M��Xr����Aؠ&�
ܝ��������\{�<<��m�kWE'Hja��y�O���.�{� '��x���G�-��k�>96�W�V�<�4 v_��T�+ě��ԗ!���'���hR7��C\��>:�̯���T'��EN����Q$���hgH=������i1��+�w�d%���\�A������S��az*��d�����Y�����R�Eӵr��l���G{���E|�����1X�{����c��⨺w-�c�t2WD�"�\h$�;mO�9�- O����m!��Mzi��%�@[�������9�0��a$�P ��l�D��q�R�e�'�~����TF�}S��T������#垪U� �)�@P� s���w�0B�,G����yN��I2��*��J Ix�ۈ�u1�Ȇ�g/-�c0��X�1��P7��Z3[���_���F�X����iMƙ�=4�"���0�����?@(#�ѼH��i��l5���ڛ|p�~�]�p��NM��=~��HN/D�8���!���!i�Q�a���]�$~��J��J����'��y��_���U��4�k��H�!��w�=���<���E��'���?h��n�~]0�K�͍5V���eP� ���8g*G����Ѥ�ۀ����fb�]�9T��k�߻_�*/ W�� ���uxMɞK�l���޷����x�s Z�r�2P�2��Vx�]Rgj�TAv��=z�A=k���@�r�Yy�w����T�
�;��=� �8ps�ЅL�9��.;&7�IEJ�/������iv����[�[왐cj((5tW�v%N��.'�V7!���\Z:���-��Aݔ�-C�u0gP*��I�
5IůV��/K�{n]F��o�sjK��l�Ōt���4k2W2�ؔ0�o��S�g\��X���9o�q��>$�l���C�7�ޙ�D�%M���@X��2�|[kם��� �P�P�4���q��ř'���f�
̪ϛ	�7�mze�z���V�6 ��w+x��޷X6�Hm^/�6Tk~f36t�T�����*. �;H�
^QK'���)����D6�s�A�%Ԩ#�F�l�ʠ��N��,���*�<�K�k�Ң���ִ0��Ӭe�弊�u&8�z��35�|B퉃��Ծl{�K���Ii�ۦ�+:�!7,m�4u,%ߖ���m���;"0u�L5�-�Ne�Q�0G��ח;J�o�bvx���ۂ--7�?SlG0�:]�-����+����BWc�m�/^�Vը�D��%��H;��]����f������2c����o.:�6޷��UI���2�F¿d�U�W�C EZ�pnP�d;�sqĀ0�gtC�~�Hf���^a]O�{����-��EK!���&���΃
��/_0�	�tZ�p�J�C���Q,G���7�pi]v�*���E��V��iU�(�Ϟ���<���/	��
�-��N��,e���YY�_(�Βʮ�5.�:r&������$��/��9:�	̹1R�5�@���R��J���h���i�w
�J�(�/�I����ƼaH�`���k���vy�+.Cc\�*L���xc�Ԥ�h�g�{�d�8�< �Gz�<��T��ܨ�򼘺��J!o��������"?˕�v�*ǯ�)�9mу�#X��ũ���Ea�C����q,��p�o�DT��G��A$>�qE�>AU)�Z�yAH8�DϫS���V��ha�k˱UD+.궒ǹ@���lߐ��������sd$>NÊ��f���TiQ{͟�;>B��� ţ�=�_~��pM�yX��4�����#��� �Y��H�(ԅ��&�W
���G�7~��O��/�������d1"I����s�{Ǩ��9���Z��1Ot2���Kl���ZG+I�x��|�`
�7���N��9�&Y/V����-ȥ%���'S	նň��W��3����	'�*F�(,x3��JU*3����U����ͦ�"34��AU�I����]�RO�-��pd
	I-���:�8sp}�E����<q�Ai����4g"Ķ���+�"�Ə�rH��-Yh��S�>	������rn����Z�v�FU��B�Ψ1���%t�J�>����<�	�«�ʓ���2\eq�gF|�{l\F�� `m� ��Gew�F9��� sN���8�CϾ���]�p�jZp�Fz�ս��'`v��U�{��X}�q�6�s��vw���r��5T:x8��vl��9W���8%�^Ȳ��-ˈ*�q��F�=�fQ��!�-J�Ԁ�.�@��K3���n�".ǌh���r� ��J�l�����QΫ;�T�����g�wwC���'3���vp�3���7�sFtZ�=I[�X���1!f��*Cy|�;m�=M�z�6 5�÷Z��m�0��3c��;�7sJ�9��p:<(
��yŃ�[!�[�9!2~>���^�r!U.X=�g���Ϗ��}m�Йz�i<��ϔ1�����b9%�w�)��iH���eh�\9x��R8<���!ke�yp�+�y��^u8��Fۼ㫗�{�:j<�uh�*Z%�td��E�̻�F|�N�X����|�hR��D�kU�'V���P`���i��hb(1,�p.���� S�c%P4��)����$lMP��G�C�P�6S�*���*7��e��v@� Oϡ�����Y��1{i�r����ZU��љ��Wl>��ⷹ�vOqJ?��d[��\�'T�����1y>t��&\@���	��-��9(d}Q�G��~~��;>{�9RkÑ{���Ws����[pJ%w��JCH�����k/77��m־{3���T�,�� ��>y���?��Q=�EwtPR�'��f�#�K���%�W�i��YKi4������H�Fa��_v{7.} 簎o,/��&J�1ځ�� ��M��%�
2� ���7ʎS��u��ǽ�,��Ve��ʤ����L�(hp�*VR�+�:]���Î��`,la���g�=s�;���dG=�_i�%��f�x��v�Rݿ[-]���6��������=9�n$�L�G�yˢ����XH`�Jh[�P��R�H�����pڐhn��O|S�;hgB׹�ó���Vu$v���K�i��u�V�HfM�I�E��B)l�S)�\�N*�ֈ���n��?�	�/i���R�Ѻ*�_�.��_i��7��dJ)i��h�2l�	"��KV������ǐO�*{"�Q��� ��e���m��/G(��/��,�S�V��^rJt��֔@�X�*�QV���~��e]Su��D���n�1�?ꂂo#�0�cO>B!�1���[<�����].��-�
lC^�.�������i���]DI������g\]p@]��i�o�u�$3;<,������=�P���{G��
'�.J��}���ͯ��=� �k'�� �ˀOl�F�j � Egā��K�d[onP`��I�F�Y��JΈ!3<�eF��O�Ax]yv|�߆8TJE
�%�Dh��r�����\�CB�h�E@�������0�6Хܴ�>���:"h�Ц�!�ba�2c2��L����j+\�{8O� ������*��_���p�
����~��l��|	�p:��r��NR��W��8ϱ
w��6C��AH�N�����x��f엸Ā_P]a�v��bF��2u@N��z���~�&�}�(r�ij[�[�����9(��E-����ܚ(��\��2?�����?�ea�T�d�K��u�[�w�ǈu�荤��D�m҆��:�M�s>s�O�H����6��h��5��p��g���l�?�5�C�Ԕ��� ����ى�"��Rh�!��5��3%��K��La��"�*Hx䜹��9;�(
�~��a�N�8R>b&�U�ES|S鷮	l�<�d���?]$�Q ����p�7!3y��*���%�,��L~Z	��Ԭ!*j6��?%�n�)�(�L��Q�� )�lJ|�E�H���!�wMU�u�ZK����\�/���I���C�AfI	
�S�ӧ��έ���Ţ�@��lxL?}�U1$ͩEϵ9���x\�2��_��c��� Y�W3�(�jk��2{��+"�1}�wv�Tj�G�*�g�h����H2�I�,��}$[�DsN2����06k��ӐNQ Ƶ���S��[��31_fN�eǣ�)�8a���ӡ0���oF(��p���b�7�e�L�~&p�Q[ڳ�6a��7�շj[!d�du�:�kF����^��w�J�B����x�"�8�1�3	N����@i:�Xw�����I{e�R�]j�P��7v5���о��{���T�<mh�D  �M��T|�uT�L��)ʹ =�i�e� �A{aw��:ڳK^�_,p�g�����8uv�1���<++�A�v��sv�!?���\�)C�.�T!�D}��*����e�(����:���E$
.߈&��(����o�h*�ix���*����@o�E���>Z��DY�w}F�\�����C��4G�%�����qJ07�?��ԧ��1��5��#�'|λ*&�S�_���'S�XÂNj�9P�08�;����m��Wڄ�bd%`$[E���D��@�=�z�&3e��]����z�P����7 �?��BC[y[�k"��c�6��Gagf�@�^3@���L
��>�?󽱸
W�pd0"���Қ门j&;J4��o�&wS
�E�/�
ױ�DL�1� �_ϯ�XX$�`��HV!x^���<v�NI�i)��-�K�*7_CHJ/6��d+�ضr�A��~����&-��`..� D2h�MEԫgY�L��������jr��E�;�j�@��FN=1h�c��Uo� �؁�:knd>?�9�������VNU�<C3���k	�y�;x��J
�)_B1y%Q_�7�h������џo�A'S�b�ǳr�t��]&��lG����"�R�9g�ܿ1��E]��i�d�H�r�b�xD�[=d{��%��_��xMfG���'͍ �0�״���&�b�Oh�L�g8�o�dp��w�8!�����r�>l��͒��6pl`�q����
���� l���a�� `�Ab)ʔG?a�������+��<0��O.4x:V����	�!���5a�b=F��prxjrϵ����Xvߧ{/��3�e/�VA>߸̪�$�6@t;r�ܝE�Ƃdn��x�������v7h�]�f?v�kb��M"juk�"e|~�u�Z�6�e��KVP��'��/�� H;b�0�kK�ֈ[�gb�ށ��a��X-��TG�4�F	��5����6u�#�6;M���r��RW�v��Ib�]�s:j7<��"Wo��YzH���Su��Kh�}u�^�,D�,�8;�4�p���ϔ�ا�^�s�cԤ`F�`����zo�%�J㩥�{0"�VvFbg�m0_9:�f)�%4^�dSx-L �$��N�]k��ظ�[�X�B��S+O*%����T���9��T.ZV��"�^' bKM��q}���`\>9PU{ާ���id�X�(U/@e��h�����,]��_ >:� �or����P7!����|�Pߐ���+S[ vzA�5e���9N�<j FF ��d�ɯ�iO���v�.�����ބ�����8NGiL�	�|�߈��]`&��!!�.��	�Dp擠nvQ�E��쨔&3'%��������۟N�7$P���a�����q�>W���j3Ҏ]�h�u����F�2]����J���全?�>:?�J�91��_
���!z��;r�0n��G@3���]n�u�u+t�Ƌ�	��9sHٹ�pu85��"I3�ֆ{\ưZ���0`�HR���:Tx;w�-�^N.D�rW|}h�W��\���h�w8���7����8�� ��
��.^E��U�|b�{S~�mJw�<�����b��ǫt�-3���R9g@����и�d4U@@��/B|�Ш��Nf+��	�����X�5�VnWE�9�>��kz���^�xR���r1�{���TQ�H���s�UBw-2	9�4��I�ZvK�;<<Yj,+|1�soiM�v�>��+�����
����'�ĂP��E������{G�@ܞ�s����πQ|R;<H��ML�'!�T�M��I��୨�@�"���]�����*���q&�@�C��W�?�ڲq��1�������n(�E���#���l0I7��Lx�"x^��#R)�kY�f��w��J�j�y�/ܛ�[n%�����`PT���\
�9�?�E����@�����˰J�1>0��ĺ-K��
�T���lv~�-2�%ԕ]%�n}9<AMV%c�`��D�X�P���=ou菉�$&�J�<�xgg�X�{��v�D��8������۶'�g�͡"�pΈ���w_��j@ϺV	"��©�W/�0�BR�~
-usbaϞ��(�lĒS4�\`e��,,]� ��	��>� doIV�Dy���Lw\�F(��ʗ�%��q!-��f�#����J�ĽB�I�Zo\ݭ����,#� ����H!&�y}��45�+��ݎ}~�=\��U��1�ġ��bF��@o�!�?���������ɏ�vɝ�n����(>�2�Dhq�k�ʰC/Y�c-��/:rl?JD��h�?�uJ���ُ�7��K�����[lK!#!�Y�eS�)����u�Ŏ��W� ���9�����3|��O��R�+��	� �Ξ�Z�bT}ui�e�e%�^vv��룁֫aD ^)I����R�
�j��k��tSN�<x��i笄]���V���ƍr2��(Z*��"�&5)D�˅pp�;T�"Qׄ
VYl�6��QR�W�B�>�S�]��N�m�/rw�X��8|�8��Fߚ!�&K8
��jr��֪�>ឈ�#Wsw����%�1|Tz�?�
�I�Òql����d��yX�d+�Cu@.��n�H�� ���Xנz�P�q���(�d>F�e�Wʰ<��)���P�P��!��A0SC�X��;���^|�s�B��y�юII_�Se�qU�2�|�Cg�د4����u�=�/�p�+nHK�/`.�X���8��T=�}�١ �dzM[?���W�K�ڕ�H�Ф�k��*�y�`�w�R�Y�J��~u�~��'yPv~�(1�ML��wX�e*��^�ç[�2��L[�h���˺�'�\��t4-��-3(=��2�s�'q�����r�œ�ʷ��k���Qy�k?�ޯ�i%o3�g������u7���rZ�߿��h��+=2���)��"z�d����	�{��E�g��$ΐ$�V(�o4K�c�`�U�ӧ��x�P�Z���9�����{�A�*Rd�k��i���B����"vE��?���ɺQƔ���u��~j�!�z2M~wvp�(5 ����kZ�QѶk�l��Nl� ��ЙrB��w�R��Y��P�jM(+��y���U����	����J�J��(a#l0�/9M�{�M���ת=��50ؼ�Ǵ�1�|�h"!׿_�ޗoW�ƻ��MԖ�*�(o��i���Z2gCut�cE�ح�硐��I�,�7$��|=�[��'*"aZ&���=��=4R�	C����'�`�~��h��9�V���3�?k�;���Mv>>�\�h�~(����{�w�2� ��/�q�bYߑE�%��,� ��w�ቮL���M+�Cmڡe�r_˞ ���3�Ǽ��%^V�G}���K! ��=[�t���[+�e[XZ�mh�+=��K�}rV�A��Y��gl��Q*[ZБ"�Y�!	�3���t+�ZI-��q�����TC� [:���٭�Tszc�%���	P�ҏ���k�A��8�����A홼6�������G=Y�/o�vsfKG�c&�n���`L��MR�·���l�_�w�����d�����A��+>����)������l.:��d�X����J�N�a'Iu�A�qf^��{�Y͓N%-C#0bֻ�����:��Uk�w�e��)�������!) �˾���wE��S|�y��FkO�at��=<wz�k�� �-���{�Ҕ�J�� ��}�	��K"�%K��d�c���ͼ��	�}�,���P��ʰ��W���o��w�<����N�HJ눜H���x��;�J��,��2�k!����I_�$g��>�~���;��;��
�� :�o�i�T!ߔ<����u�v�t%V�f�I��b�����K/���+m&o�b��ԯ� �D��!�G^�M5�8�u�)�Ǹ��Asw�	����v	�H�V�<NQ��l�㥜Ԡ����L���w �J��1؁B)��&�~�.�!�v�8����=���P����˧�Tڅ�,Je�7'S��?Qe�T-�j*��5�,�O���+	�>'�D� E�����k���(x�m#ԝ8�1�@Ή�\�_D���/���R�8;.��q'����6�� ��W�O�\�E���c�)���Po��4���;�]j�s	�9�	��h�N0�W���xT�����"��T`�Ŭ�
��XɄ��8�����g�p,��^�����h_��h$�~��X?Y&�`�W@�g��=a���H	ϡ�-�ɰ�����݊ӵdpGPQ.u�#QLu�U?"�ËC�!F��;�M� Uا�v3"K�<i���j</>�%��@4�˝�n�q��C�U�b
�g�Tc��U��bJ�T%P���d���!uD>�'����0�ae`�(����E;[��8��Q�;�|�ک����| E'���xG2�Ǡ�6��_��t���`nYa��m�r]��:���eP�O�U\ꅏ��伍t����f;hJ�ֻ��z8��!~e� �cR��D��>(�4݆�]�S�y��n��Hy��;�E�d�I� ��r������#mW��1G}�gHB��l�)�4��nn�8��Nr����}$g�!z��?�⍜�$�,sbQ� zہ��-��F��G<�*�a�&1^X�� �:��_��UT���|�M��"�t�>���PaB��SbT�Z;걯ao�0�T���7aa��q�W��T�W;� )��t����%�:�7�J2�闡1�%�zX��*�9Y�=�����z���M�� ��YP�M�K��=��t�Ӕ�ɋ
�h�y {����)6�Hj�4x8n��s��Sm�3V_;P��T�LX=���'�ה�4p�����g�3��%����|�|��b�&����IVxk8�@R�Wj(a���b���J!������MǙ#I�$5}^�`7.���o��?b7?�]�Y��%30n��ʥ��Y>�������?�ʦ�Rz��� �䳙����_jL�h|�X�����E/�.���^��II\�����34�j��@ �^@&���9���~_ �?��3}텅#3���9�HK�x�YZVB����@��6��r����?�l�n�r'镑-��Fd����|`^=hU��i.�]rX���dH��n� ih*���h��\���8fk����o}Ƚ<�y���4�lE.g�9�3�p��4_Ɵv�_�h�;*��jm�Crq8�f�v�!��:���W��V���[a��`�<x#EZ��-��Be��~��X:�I x�����!(p��PVLʚ-{}�i>m$j+�����1m�	�֞
:�he��j2���1v^"o0D�$A�` �\�_�U��!��c��#�&������c�k~�\���uX҃�;��R�.��Q.�b�00n�	md 1�hAͭ����Ն3�/�G�>5BϪ�I�4."�+C%ȶZ��0�rx8�	5%'�?4a�����o�l�g��p����eu��f:�*�`}A�m�NI-b�Ⱦ�pW dt��CC�]4bWa�K7�~)}J�݊xZ�i�[�a��i��>������ꌁCsD�^��qq��(�o���9��kM�C�4O�3�d�I�I���AF�k�_]�y=�"�g����#��G4UHtհ�\H6����.�ۧ�t�eRV��~R�qT���0�Ҟ��C�6��~
+Mh�ϓ�;���~���gZۗ��L�#�R΢�uU�`M>潷��v1�HlYt�l#����w�Q�R� �p��m$D� K)壞���k��*�I�ː؈�'���Z��1&R������z�ܽ5�P��j��ux֖�ϋ��q$z�/dVe�H�0�t^��>�L�BS�vX�(j��;E�z���t��B&��l��az3 9��;���{�.������N2�x��, �z��Չ�
�Q�\Wҭ���#f��V7+Fz�=��52*�p�'�#�Q/��=��aY5����i�Vt6/-J)��m�VqΘ���桫1������Α�~m�UT�3�d,������j��_�犏�t�ZB����q�?`!w�V:����n�ٷN�>s� ��E�	oϚ��ZG(��)�\QӾ��<0�6'_�Hۭ,�4P�&�Dy:9cP�Ѱڷm�x"�L�W(��K�i���:��<��j�Y`��Ų͇��,��X�A�nɣqG	��/�"�2i�.r�p�(�w�1��Y�5���L7�8F����Wu�����ҏ��ԱK�y���0�]�	GD4��d��Vw�S�ʔ�8Ʌ�Phy����������[��.��� ����w_�(dΓ��u󓩭 H�^�[�+�gɕ��D�J�q�$�K��Gu5a�2}�s��;��'^9�=Nf3����3���ȗ������G"�N�o����
�Gsu����(��K�e�r����4�u9� j��'Y��q��P�Z��J O�m3~5\i��aU� �A �b�}L�Gfw���J?Dm��iL����DVO�ֆ�C�DW�qva�9��K���￱4&P�l7o��jK���WS�,�01�5Hq�3�,a�)������O�������� ��
7�D�i��� �$+O&�� B��ɢ��I�	1Ǔ�Q��1�H��qdh�������,����P�>���k��{*��b�Æ��q�����YR߆T3\��H�ĉ���f�"Y����k��o�R����KQ�bֵ�M��By��1��&�u�<aӍJLXB'��>�����E��`�>�FK���"�~�o�Ͱ�k(�(���Q��ԗy�(h�}6���b`��ل�jW���T�.�nXց0Ϳ��7k hTX5~���H��,�6sF�O�ez���¨*X�,JRjL>�����k�)p��g�U�s25|-�֧�x��ǹc~����ҞFF���9����%�4˚���GɿqRF�)�웝5���;�Υ2Q���^מ��l�{��u�7)�v��+����=�V{.ТpKL��s��w��g;�|o2=W�*c�4������%k��ߺ���a��XD@�X��N�&b��"���3�wZ���\�n��+�*�V\��ZqH�Q����ʢ���L&�{`!�g���8���t懥]���P�����+R�J�xҮ!R��c#����8 ��w�����ދm�@��3\~}����vi�5���u	ᆠ�+ט�괔�'��i��v��3gn>I*�l����V`�嵖��{a���>9��n���u\�#���s�5����g���AVr��`����|�,�0��:�����~�8$�#[�����\�G�Ղ�vkA|�px)��&�L�e�~��]�H�C|1g�>�.D~�hU+��X��1R���o:�SFN*�cp��l۲[�;>�)�7�þ��{hQ���B"�AJ�%��k�������쉿�!�͏:�+����3n0���K.8�<㺕gʱA��Y,�;��}8��Fʭ��}��$q����`إ._N��l�Ǯ�%�޳�`�*��5�n�Q�7U�R\믁�){�Q�˗O# ��Q�#�v�-z�[�	JH���v��=���R�L#d̯TjJ3�>�1+y�C�m�%`�݋D~v�C����	������!<��0�u��4}�3:Y�N�%� �N�EgS� �y���vc]D���� ���j-{^��*h�d��`u5jؚ�����l!S@�BG�v�'���H/R�������רp:�E�^O���;���{�=��3_���3�ʷ�=h�t�;�0nB�� K�1�"!<���ũ���j6M�[��F��yVw����x��������Ǥ�w���^��MOk�1`�1}�R��N��|�CV�;3~Gw�����H�~�����|�3�L,)�u�#�3I�p~�~(�~C�Қa^T�X�[&ˬ�@;_�
<9\�q>a��o�I��W���q�Sc�D[�h�*́4�����q�{~hkD���d2.�|5q��1��0�GY)X��ҟkBqs5N�h��Xxİ�<�g�W��`�<A������<��UGe�S��3,��P~9�+�-3���U�$�Ҩ�(/��-?V��E�c.]��U�v�V�NyV(�a��^��s��xBr��]rbbe�c�V�Dၷ�Z$�������YM��Js�Ԩ�\�{���@O��1�|��`E�y����{x�Ʈ�%ie��rZ�e�)H3%Y=&2����tĔz(��yE�JV���Ի�`saK�����-���s�ɹST)B<l�e�mSyBv�����߽�}Ҹ�"�Ğv��?�i��z�[�d�?tr����'���t�����e��EM����7k��q�<�W͙�$'-Ei�*��ߕ�_-aڳ���<���u���|,((�V'"�#�NB��W�	:�}ڽ	w��k���'|@`cy	��'�� ���ku������Nۓ��r]GM���YC�JIK�\�_K?u���r�����"-:?5�[��%�hK�?����p`�`3z�ڨ�\`��O�o��t`�2~��X;=?-N��n���w���_���>fob���o����C2j���9m�g�Tqї48-�H��z�q�P�Y�t��a��k�����ж���k�N���\���P�j'�?�c#��޳ �]�p��%/�o�i�-=ڢ[�DXG�,Je� .�������}��i�,�~��J�{���_���|u���<����HVj8�T�]�Dq@�5�	�p?bC�qȿsRd�
�뤒�U�xf ˫�+���)iE��Yu:��Sf��.��5&W\��a����" ���[�|HD[�t�SJ���
���'U�'�/<�����5]~�?�zm���:�p|e��$��#r}/��.11l�H�k�y=B�S���j�����&q"Dg��]��Y�T�B��?8�D�	����d��T�~�»� e�����H �q\�>���&/BB|A����sDMEn�?��6����Ja2JQ�s،u��`/��p�(���,,��^�
� Bi����[Z�8r�N�΃d��CH����Dfvx_X�5)�J1���e��SJZeq�Ffa+bem&Q�Ђ�y�`�$�SE\2��1��%ΖT
�ˌ�6��gٚN���S���r��'�3˹��Sd8�x�i_Q�RB+���^ +�u�7Z4��餓AJ� �q,B��u����1f`� ��a�x���)��o�1�)��P<}�`����ҝ�hk�U�ۼ0���_O���,����j5���e�ܫ������K�㦏�8���d��m_z�To�AӦ�sL ��0"^*+�J���kF�����B�����LM�� �}	��R}7PquWw'mO���:�U�����Y�xVt��+�`�PL&أ>;�&ǋ���y|l�c�����q.]8�D姃�;@����������c�v�r�׌v��Tή*��1R�ׄ`b�%7�L�y>�i[!LK�p�>?��n$k_���H��ƹ����A�\����|��TC�&BD2L��v*:�6�?��e�d#[1[1��yн�7y�qD!(���r�[|z�Zo�L<��e��N|)�OA����|��o�"��$-�����ty����sz��}\���$Zw���o�.r�=�"o��C_bI���}f����O��njf���!�O�Ov�- PEt�����UyJ���)M�1�u����r'�N̴�z�'5]\�r���\��z��W������M�w���Q�ͺ�\�DDb��S�\�>F4�s��3ٶ��g0�bZӵ7_����{���{Q������e9��0=��������*3(jp�g���N�Ơ�%.����| �-���Rs���z��k:�ڷ	`����h�o�m�BA����zǉ��b�}WL����)��&gۮ��Q�;Ҳ?[�l¡�Oq6vJ2mHS�2����p�_Sy
Ɛ�z_館u�S��t�_
��f�ϔH�"s���j&ǙHW���9m��:j��pqeL��BEV>if����R��d��"�.gB���Y��h�) K�Eろ�K���N�u��xܠ����!{������ فϗet.�V��!�b�����a�';g�_{B�Nм�nnGb�����ň�;c��-��Xܗ�c�^+.I��׶h{Q�����RwT�v6v[�J3�n~P���-��?j�4h�5P�T�uo�df0�:���v���aIX.��Xٛ�b�~+|�hn+��"%u��z�x��>�.99� �I��%��We�N}H�\g|B����"���'E�Ig?z�9v��z��?���������Xv�BW���e�'ށ�\�a)� +�r^%���O(�lX\�|�q�	��ޒ���n��n����[�Q6i�i���#��k��L��` �nw)5_�1�f��e��x���W�3�N���0�5*Իz�%x��]��)3��uџʼ��C�����Tz���ATJ�����"1�$
�I����J�ogX�ج���D/%G)���L���V��Mj�"�#{줗�1��X$��Fun��D4����:&��{O8�~����h%��<o6�X�!褈S �Ж岼��������9qP�8��2�Bq)�v��(R�~�
�j=�B�ii�
ch`_]f��؅�z�YږQ�q����g��ٳ�80$h`��ø=֌�QT��j|4#tl6�@�<�F-փ�����T?�J?���@<i�<���Fʒ�5�w�H����&B�1�򗳅Jr�y����z�\�^e��/�F�~Y�3�GV!��t����&fY"�����N��Yb&�(d���{�L֜$d�y�X�;s�djW~N�'ݏv�{��q6��� ~��<e�2[2�kL/o��|�T,][����u6�M���h!��,$L�k��c�E�#reA�� y�M��J�$H��Mh�(hC��.��!��Z�\~"�����w��Pl���t�#O�cȧ���������^�}��9��o�m�Ax�� ꭖ�F6F�&�g?�ʊ�����,��2��F(j��D���A%7�,�ΤV*u,������M�;̝G'm^-f���p���1�	cO���T4[bv&'�}gn4P���P��w0q�����p�Ht���\�}������	�&�յ%E&�]wpP�)����ڊ�L��>��_�8)s^lfjE���\4����o�{��#�u,��"�<Q�u�;{l��N����̟ɯ����#�����`��uf���+���QA�#jQai
�������m_��Oj>��e[�����g���b����̥X��V:�+@ߌp��oOɕ�,�;��U��DU�����Ō�W�Wh�A����>왯E�ު�j��i.uk^D�(S@�d^���Ü1E��.���8���lX�g�_�)��q�c�n�Oeɭ�w���ˤ�k�<��n�^�g�H���	�����ρ��N�9+��
n6��mv�*����Z���=9�i��6K��N��#�V�%lQ��gUU����������{at��X���/����z`��kU�)��M��������M���Y���: ����#���M��v&U���r�.��Z6B�Lv�L�VIt�7!���+U���K�8�����t�t�2|�".h�3��= y���J�bĻ<��������E�.��4#��pt�O�o�_�[_��m4A<�?^T~c�䶂����]G�����i���^�`q7��m����	/{�D�<�Lɤ؄��>T�:x�G����L��T��E�hv=��E�����|��r�%V�5��Ɠto �ػd�R���k�x�����ʦ�I<���d����/I���E�憠�;��~�3������z;�.;�;�ړ
a�+&������j�"�I�bI�=	���`i�n2��3�4|��ǩ���<������0OZB�H���&�#UЬP�"=sM�ɡ����6'9�d���Ӵ�2�I����h0�J�E@��TQ�&ߒݽ\��:��h<����N���k�U����tmk�d��h�sb"��v�LDl�����Xsw�'l��� d��X�2v_o �C�x �Șo]Z9��ԩ�:�&I�TĆ+�Xz2���_�!��1k�Su�bk&,C���B=V�<l$E���
�/�8�{��8�ｐ�m
<�����J�������o2�or?��~Q����U�өY�T�:��W�w�ά2�!�����5�>��1�`���R����,� ޢ��~�� |�����(=�F�I�q����Ϧ��__��(�l#�+7p����EB$�<�(��AR)�a��5�4����0�I��;�oX�禍��Cu��(|�0i:�Tdp_�1��G~��a�(���a�0Gb�BD�M����0rjL9�����'�N�X�'�rx���9�L
�. "�F*�%b05��B�M*�A��-�����k!�10���
�y� �z�������0P����8mH�h��JP�y�wܭ�Ԭ?��G��־ W\D2�N�R�Z��{�wU�-�TU�Ǌ�]�6�Շe'�v�k�-`�x�_���T����c�_�㉰v��p����H��'�ئ	���)w�茶�B	 ��^�j�9�v�s��[�A�,@�ĀI5?��YKp�M�:W&'�Ʉ��k��$+���U�_��\��ǁ����a���5x���$�Y�(f��]��]q���&:	r0��9Ze�����._�0��Ds(�QK���>-ey)!�)<������t��s���?�JV����,��D}Cw��&�џ"m���f�\$�P���y鲾|\���A�W��k���}�@�Q�X����,����l*`�j�Au�O���լ�h����t߷rxɣ��I'$�{���$���x�VemL{�n3�!����R�V J�I6��;�����;�6i�x��I�y�:����g���M��>�Dv���4j�f#��d��x{]r��(zv�c�zP���d9�������&��)���?��b�Bs<����.l��J����"ct�}t�ܺRx��޸��ۖ��{�`�t�Keɷ����x���;#׉��Ծ��5�dS�@fT�ee�Ha�(���������W��Ĩ͢�V@aъ�R�����;��_�f��q�	�*��q���3�����~�������}���2� ����-zC:y����²���
�.F���O/�{_�v�iݤƆ���/�Ơ�"|�����|)�,�0V͏�}f� �A�ML�l��$�P 8ys�چ������k1���mx3B��Z�dąـ��M;e��N}7Տ�m��n*Ŧ�8t����]��*�"�_s��j3e[Ű�׸/��H��*զ�m��r��^��v[m^�^�Yh��U[PeV#�Ꙧ�A3h�0���E!Uy�C�Ьx�<Q�\#	cآvk�v�Ke�*�,��a���D���OOǽ����)���ƻ���wc��dd@g�Qn�*��!X�"!̀�44|�Eݝ�[o�٪���؊"~�
��n�R}��o|��蘒z^Izb+,S ��So-��u3���;6i'��E�>��z��� E�Y^�O����EŦ}��|�Ň3|͗Tx�Q����� X�O<��N=q+x��q��pP�iKWjaU@��t��|�	.Xou�̷|�����>�7�~R�1�JŤ�SO�Q�v.H߫ O�\���	]2F�6������k>�y��D���ŋ��5|,�B��ޢ��N�п�'��$oDG��\�?�usUH0��Z���A��j%�t#�I��y�aI�/'�R���A=J�F=��3]͌����/��ξ�"�E̳�J`��怣&�I�r�5�L��[� #R�KH5�����$�$�`1o�����Ru��jF�������zj\~��Al�P�V��=8`���x�`���;��UX����H��?��js��)U�m��J��e�+7�u�z�M�\�x�uq�`�L����xBs�ix�%܏��hDt�d�Hn�?���v�۶K�UkJzѨ4��ޡ�M���!���ݪ����Mɦ&�X���,`M��B���LӢ���&�>�vMnq{�*�����-,�ak�S��k�U�o֕~�8�HQX\a��ɢ�F2�l��C�m�E�t��5�3�����KD��z�z�U����"��:p�Ow��}���M�����S��o���p_��}{�L{�:C2�$Mt�Z��B�A{'YT.+F���� �l�"���	���Z�^���[,���;Y��#7�j���e~�Q�l-��!�zl�[}���؄\&��H�b6��K&�(_�9M#�n:!���YJ�wS|�i��&�m�3j�L� =�6����џ�r�i��N
��5�~\�O��#�j��.�Dw����T�kasjiw?�D�=WY|kK�y54��~�"�����>!�4Zǵt]�=�4%T�0dM!���s��FXrc��*J&�i����=Ņ��s*E�؉��6l���Y�ӱ�2��m�7���[J�7D�?A��dy	���(6���͒&q}�}�,h��I�b��I��Jz{��p]����-[U �؍V���}9����U6�M��|o�U��L��TY�8{�CT�ג���H�|�
l4�Ӑ=4xQ�jR)�Β�^
�x6���>`��b:< ���ҩ�������P��ϛ�tW��[ݼ�z�������)'��PlM�,Wf֛�;�eFS`X�{��ٜ'����u�3����+�?˴�n�Xs��ə��$�D�m-Y��-�����f��'	���K��n<H���Z�	�ރ� i�?�����a ��[޳iqRѰCLyo�- ��~rA����LuU,s�	g~���Ԍm����>��W�Ʒ�r�0=�z��ν����[ʴ���6\+��Puw�j��~=9���>�-6eU���1���Cu`GQx�?�ֶ{&�U ӕU�=��iAzeNf-�t1�#��R��D<�`0���	��FM�6���4�7���Zbs�AO#r�܊�6'7��|s8�� ��m78�PUK]�k��\��Yփ�=2�.�l�scE˶�m՟l��Ι�2�vՇ�k�j{I_�����{xꝰ�N��A0~�h��=~�LZ���}q��,mƷ�ed:l��2����|S�e����7`��>
{�M��!Z.�Fm%S}�&��>��I41�BE1h�լ�	�En���t\W�^�d�5�������9j��G@���Zͦ��Bqa�2��^O�:f}օw�S�(�􋏏�s6T:�U�\Y�a-��D���@���rQ�BZ���URN�c��h~�{�P��$�^�S���B��~G��̐�<��Kf8�m�+�n%o����G��%ۊ r� 쭧DH��&
@��]U���_�T)B���e���'� <x^GPH��q��hhۅ���ʰ�v,�}'�%򇧓E�^�����=�vL��o#ͬ���@��ؿB�[;��SϽ���Ӯm�
��y+r�'e�.�k'xŘ�vH�l��Pl*�z��QZ��Ez�����X�լ��}����Q�y���Y���}�"��E['P{�;��m7[�!��:�U4>���;��dsv�m�H�h�Q�e}޾�?\l1���Nc��ǃ�S���^]E���f�3a�f=�2(?���W7MH�8�"�8P,[~4U�ާF�Wdn�҇ߓ��<}S[�}�mZ��Q�߀��4Y��h,��$r\j4KXcLB�0_�H_L�p�v���6�nёV����~4����/[2������A��=�n���{��{�|9��j�4e7��^�F+"|5�����so͉1��ƍ*���d(���b�FA�k����&Q �����Z	�pR/��l���`���a7�m�$��IzK,d��r��sT@�{F�Vy�Hh��b�f*z��솉�-ST�,����:��LtC�M��)r��r�{�te0��L"�XGVD�W�� ^���@��X���{O�Ϭ�ڋ6ґ}����-֠|�u����t�&[���h2uϙJ�2@I;����)�ָ��d��wU~ڜ�����+�u:.�M`PI-�����V5�kK�Poж[�}v�\�6.�'<@7%)Ly��Զ�Ő�-BY��Np���#v��T`�ܠ��� }t��4r�Ȋ.2��#����\QL�]Ʈ�����Fr�����e��o�_�b[���]�F�p���� ��H��x5��	}���M|��t9/J����Y+x{g#�����:�R�8gL|��ҧE��%�R�W*������% ��B��D�B����$kBW�@D�����]���(�8~� ��O̦��/P�Z�������1q��+w�Zx/��p�V�_��;Z�$���B�7�	�Ţ��a*0y�n��E��<�KXӛE��ܾ���E�`����Q�8"��2����X�����+�m8�*W�5���E���E���0A�^Jܪ���ҚI�J?�I>�����\k�>� +-���:�;@���5 #<��#ó$i5_vY_m��t�7��[P[c��'>��Y��X�Y|�<�P2N�0�0�
I#=��jR��r�W-F ��M*�b�� �9�>|�]\��OhԷ`����~,����H���z�ZbI���Q:�}�)-m& S����R���br6�KHɠ�7�Q䑧��l�&�<��&a3<�k����DCW�ǥp�X�K�>���H|�bG��h�_�,�{EcTn~��O�\m�U��Jte�}��e)j&*f�Bԛ4�6��4�W!-Z�cZ���M��\t�V&n���Uv�!�-��ur��'��ꐷp�>'9ZS�T�<����)�qh���b�D��U�ϖ�)m��8N�D����P���H�(=1Q�=2��^���mQ�?�%��y��i�j��#�/yK��A��#Flt��0Dh=�J5#��Y�qhW����c�lw�N�S�E��9��BW2�!�ɋh��R���b�������Ժ^���Z��!/' ��KƉS� ��`�I�z��b~r~�eC�Z�
oq�D򢳞)��n��p�8�������R��l�<p�l��$��?�ݝ�ߪ[��N�M��D�|1���d���J��x�\u�}�����<ڈԒ�����A�.R���
>����g�ф�D�`H9���@��:Y�=S��t���$�ʶk���)���d�����h0�����X�<tͦ�Bt',c�t!��ǞB[腣�N��Y0|�Z�}t��<r�:dHs��ӥ��.5��m��T��aÞ-�U�:=-��
|./%�Є�X�[f�aZP��F��OW�Ț<XS�M�ʋ;tTZu��N301&&y@s<�k���붓��ϯa���E+DT����| ��p��ڌ7LeZR7b�C��K�`u�OʹQ��������g�@{�, ��Mf�Y誇S���..��?���U^#�Q	�X�6!;%�R�N�V)�Q'�2kC�