lvdsrx_inst : lvdsrx PORT MAP (
		pll_areset	 => pll_areset_sig,
		rx_channel_data_align	 => rx_channel_data_align_sig,
		rx_in	 => rx_in_sig,
		rx_inclock	 => rx_inclock_sig,
		rx_out	 => rx_out_sig,
		rx_outclock	 => rx_outclock_sig
	);
